// Verilog netlist created by TD v5.0.27252
// Tue Feb  1 03:21:56 2022

`timescale 1ns / 1ps
module ip_rom  // ip_rom.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // ip_rom.v(18)
  input clka;  // ip_rom.v(19)
  input rsta;  // ip_rom.v(20)
  output [7:0] doa;  // ip_rom.v(16)


  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hB0D6A13C038D1FA7BE4FBCF7D55153F470B627EBCEA6D49767FFE9FFBBF9F9B7),
    .INIT_01(256'h3239AB1DD37DC9C96B8A7D655A6C9A247F6EFC8C5E36474495B745D25AF13BA3),
    .INIT_02(256'h442CCDF56A2F76B0CDCB7ED323184443D0A37714F9C1E31D2D256A9148B5DAD6),
    .INIT_03(256'h248A31E2CB37E1FF6B799D2A5C1C44BA249001D6254F661912225A4356E52766),
    .INIT_04(256'h56A75AA4DD5E95F1E37DDFF87A0F35730F7BAFFEA68AFE91820EAF4B29A48E49),
    .INIT_05(256'hB382C14B0BFDFB69B83AFA8CDB5A5FFC418B2871C0CAC86EF4DC1AED9E0D5BE8),
    .INIT_06(256'h559C120281E47AD70C2CBB5443FCB3A10A4084A85520A54AC4B28EC962291553),
    .INIT_07(256'h932C51BCC9BAE69E5CEBCD997F0695EAA569EBD2DD8DBB5DB630F4E68ABEEF88),
    .INIT_08(256'h425F26B160F5A8B156476C0D6E02295555F667F0BA203AB9EB0B7554BA863DDF),
    .INIT_09(256'hCF84541AD74AA8363190DADFCAF6AFEF158E764FE733E173BF27ECEE66C7E4C2),
    .INIT_0A(256'h90CC6879A9025663B513D6309139CE17B40B1539827CF73E64EAB49A5F43ECC4),
    .INIT_0B(256'hF86E43623BA3A659064EE5B4DD1B5DD8006FBD84AC54BC92D8D3B3BC64116740),
    .INIT_0C(256'hE69A520876F6936C44B435AA1BF7379EF5C0D53CAA1469568FC55CC7E13CFB3B),
    .INIT_0D(256'h112EB7FEEFE9332BE623676F9DB381221AC6108C308F218B9A9B770BEB8A10A2),
    .INIT_0E(256'h59C06C7C009A74C31E65499DCDDB61CCEB3343D9EB18EB7FB41A1CE60F77F6F6),
    .INIT_0F(256'h9F7BE3D73BB92C4D656A9B67DB78BAF0BF7EBEF3DF33ADFF8F97FDFD25CF76EF),
    .INIT_10(256'h7DDDCE67FBB769557F7BC76EB93E9AF0C913CAA544F77C5F71F55ADFE986779D),
    .INIT_11(256'h7DCBB89A983747E47DCADF51267D84362C2FF44669A3BFB77F5BDE7B6DD0B635),
    .INIT_12(256'h7A8E61C6A789C55BF9272E750E8FF7EBD968EA7FEB7A72558B0F3C62F61F74F0),
    .INIT_13(256'hD9C72592C1FDEFCF57C33AE3EE87FB672B2EF3BCDFD0BF658FBF86D2E79C3730),
    .INIT_14(256'h71001E21A0A8C5F7900C5F6D9D4F8218EFDADDD0589F65DACEC93DE4CB6603E5),
    .INIT_15(256'h868764BEF1DF7DE773B7FD867483CB724DEFD674DAC9114C7DF77B9607DF7BF6),
    .INIT_16(256'hBC7D57F5AFF7B8E264690CECC253022479F7446588AED511BF7ADDC0878FD294),
    .INIT_17(256'hEED71B91E3E07DEB01FCF5B6667911CF94C2E5F02E254DFE6263FAE9B15FFFDE),
    .INIT_18(256'h84CAD2042ABB763B9AA78322DF20075D1F69F8FBFEB8C83BACFFFC7CE5FECBFB),
    .INIT_19(256'hF19F9FB88F000A074FEDFD7E0382775FEEA6EDFFF8DD6661CD7B202502BFCFE8),
    .INIT_1A(256'hBBDBE6CC2C7D6ADAC952DBFBBBFDB6D647E5B51044D97ED222EFF209689B37FE),
    .INIT_1B(256'hBF8C09E417A417DFF0217C0A0B6F764ECB5BBBB3564F104D54D0DBB6EF651435),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFECC56024B3001CE87809FBFB8383935B6CCEE0A001),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_000 (
    .addra(addra),
    .clka(clka),
    .dia({open_n69,open_n70,open_n71,open_n72,open_n73,open_n74,open_n75,1'b0,open_n76}),
    .rsta(rsta),
    .doa({open_n91,open_n92,open_n93,open_n94,open_n95,open_n96,open_n97,open_n98,doa[0]}));
  // address_offset=0;data_offset=1;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h10A772AA24689A05249106C99A638C12F929B885E3C40596569A0DA099FBFBB1),
    .INIT_01(256'h7514E60DA4ECD0472A71BB5AD810201EBA3AC98AE4824BCA1505096329827E12),
    .INIT_02(256'hFF18400ACE054E9B42860DE320148A0B8AC5444978CEE4F65CEBA2E1792ACB14),
    .INIT_03(256'hC965947B945BEE2DC09BC79C132C8F1D24F001177071554606AA9272B6C131F7),
    .INIT_04(256'h57C9FBC67CFE7F83F5F9682C8C73DCAC610612004071CB47507315B0D6F234B6),
    .INIT_05(256'h3657B5B5EE284D9782A7ACE7FCE5E002967CEECF2D2EF3B3193D8332C4976FEC),
    .INIT_06(256'h7E20A1C6FA0DA9FA5DDF24BAEF09247EB7AD6ACEE3CD9BE1ABCDF5F6DDD4B2F8),
    .INIT_07(256'h4840BE0217094B32A17E56220456CD7F320ECC195BF7DFAF6FC55F0213D800BB),
    .INIT_08(256'h988398D58C92E509311CB6C0B34FACD99D4D8016E295F74BD5A013F7F67B1368),
    .INIT_09(256'hA17C71661CB2455B1D00A120991B201227F01BEDD14612144A683B0002518054),
    .INIT_0A(256'hEF21A9E5509559140B60FD55AA8921C16AC5289B57420C831B054763F8BAB819),
    .INIT_0B(256'h8BDDDF06CDE41B77DB1BDE5D6F20A72ADE8ACF69274F8566F9E560BFF833DA19),
    .INIT_0C(256'h1DF4E7610959366DE102D886F0CC84E33E70778BF9FCC23C444A7B71D58A70EA),
    .INIT_0D(256'h5891C821EA9A60D069ACD0105260F7FDE5FB4EFE8B6B943B6F264166F73B2FF2),
    .INIT_0E(256'h83AED115AB551AA87D53B30587D05FE5F7C336B61FE3F443653EE2D7C049A41A),
    .INIT_0F(256'hA30AAA4CFDA205723CFFBED9748245BBAC464184FAC64680D1E817FFAEF1C911),
    .INIT_10(256'h8662A29004DDBCFF001A8CC1F4602073DA4B1B59D858C081163EFB7F37B8DEEE),
    .INIT_11(256'h937D4B83024938CB979B33CE8D84E9CCD2C07193BBCE7E0090E0E9800665E384),
    .INIT_12(256'h9FB0BE1C3257F1FE6892D388B15548624243DE000190845FD4F2F19D9D65C77F),
    .INIT_13(256'h137141828A43434BA6ADCFE62D99A64D5C4DD4CF2405F009D7CD692FCC06FC06),
    .INIT_14(256'hF9102CF501C183B836A9372BFF484A5304E12652B2A0CF249891A44E106C4A75),
    .INIT_15(256'h9BB0804584DFE688B4F81100DB28204400412080841CA6381DFE34ADAA6D7C2F),
    .INIT_16(256'h5E87F858795A6B486D4060F692053A84AC78DA6878F03E779BF9831FA83F9EF7),
    .INIT_17(256'h1061C0F173F30877E47C7FCAABDA4004B22C2712A467A1F0EEAA61444B3F7FE9),
    .INIT_18(256'hF6A7A5B2E449947DFED06D7920E291A4040341E89305AD8459CA2DFD9A709412),
    .INIT_19(256'h0EE041400FE5BE218251004977548C20010134C30E60EDB4328C042480DD80EE),
    .INIT_1A(256'h4C34B8CAF419D0B460F8323444D22C0897F521BC1DEC4F097119F79655424C00),
    .INIT_1B(256'hA08040AF7FAF7DA7D487B52C3440F49891E2132474D41D5488B6E610103A6086),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFF7102D2595C9703C22C0B4F9AF8788A20703ABCC97),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_001 (
    .addra(addra),
    .clka(clka),
    .dia({open_n130,open_n131,open_n132,open_n133,open_n134,open_n135,open_n136,1'b0,open_n137}),
    .rsta(rsta),
    .doa({open_n152,open_n153,open_n154,open_n155,open_n156,open_n157,open_n158,open_n159,doa[1]}));
  // address_offset=0;data_offset=2;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0284B98003A601538298ADA995459704FAC127CA495095248554115F08F8FA84),
    .INIT_01(256'hEC6B376A6F175E7FEDAE5DAB7FABA5B7D5C5553442500B87983855F740F1E882),
    .INIT_02(256'hBB9DF14AC2988902AA88832FADD3F9502D7D3B6B11F82548DBBB4DF43C7E2C69),
    .INIT_03(256'h4B214C47DC55079202E00A948414849C004053067740626106AE84A3E979CFDE),
    .INIT_04(256'h974FA1710331A87D2402030300DC0362D763A367B7A8C4115F5F02BBF7E88E92),
    .INIT_05(256'h8913CC47300199C638B258FD3F39FD59E73E62638D623BF0C01D02241C200161),
    .INIT_06(256'h79505BA2A384522939F3C0DA8C0577C6338EC6B661EE89E8AA3F3B3E3F383002),
    .INIT_07(256'h7BAC2C1AEEF094A23A956104E23414448501C302C93FBA2FB3E5AAE6C15F4288),
    .INIT_08(256'h2F5A9895494091C48044043C3043A4CC8D000B200EA4CD23AC2A60A54A982A17),
    .INIT_09(256'h6A087144B42C13CF4C2F38B370C50AE8441C045A267D0567106805C66111E065),
    .INIT_0A(256'hF7E948076D8AD084911E08E119320D7E50FA6522AFA3CE6CD5D274B8A45783C7),
    .INIT_0B(256'h368C277222C8FF90BD750623164FBA9016E105064D7432F708145B1586109F50),
    .INIT_0C(256'hC297397D12A5A5CC7EB5C00128FAEF5D831428B254EB59DC2C3308062F33AB54),
    .INIT_0D(256'hCDB94B961507DB13E96034FEBE5B35C4339CE394B3864D8E15399E22A08B6328),
    .INIT_0E(256'h11CE6874678E78731A31E69A1D9FEEE7B0B520A9D4B8ECF3787A3085907E07F8),
    .INIT_0F(256'h917020400304511D944538EE456A0967D03C200802748432968FA40CA29C165C),
    .INIT_10(256'h40444D5EAA80760AF6C07ABD4D5D36B11046826D4011007173CABA00112E9101),
    .INIT_11(256'hE401720A80AB8800E782B47F3ACA697E109306822EE4034C3BA730C9FBE1D998),
    .INIT_12(256'hE52023888C3807A41424A44678FA8600318334C702E0E34A5A5C0182AAB901CA),
    .INIT_13(256'hAEA674545722829D735E5D38899E05BA1EB302608DE548E81D605CA511A63344),
    .INIT_14(256'hAE5574DF46D6E9B258AE967AAB7575AE1AD93BB8D4B8BA8176EA31946B9A9520),
    .INIT_15(256'h771CE2741BDB601737A8E70102AE006E039F59F5152F14206DB677222ADB7D2A),
    .INIT_16(256'h2582A80014840B0FA9507AF0ACAFCABB2F375C6AEB6570119B6EE104AF8F1425),
    .INIT_17(256'h5E392FD4EEE875EE61FFB3BA6308403D3E0D083BFA6F6DF088886907ED3F4FE1),
    .INIT_18(256'h1FE16174C220EA0CCDD7DE58AB7088BFF3BAD2F80FE969F5158575DB1FE0D7F3),
    .INIT_19(256'h8D7ADF700F891EE4011EC5FB17C5503D2FC806F3E2EF450728E60084801EB042),
    .INIT_1A(256'hF71F2EABEC121DD7FF5FD53FA783F08082B97F4E99E5EE115AB5D7954974FABE),
    .INIT_1B(256'h30AD282E3FAE3C2580A44023257C0776EAAB28BA4B3413B573AC406BA802B9F0),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFEB914101454E41C5F33804B2A8500AABF31C29E4C4),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_002 (
    .addra(addra),
    .clka(clka),
    .dia({open_n191,open_n192,open_n193,open_n194,open_n195,open_n196,open_n197,1'b0,open_n198}),
    .rsta(rsta),
    .doa({open_n213,open_n214,open_n215,open_n216,open_n217,open_n218,open_n219,open_n220,doa[2]}));
  // address_offset=0;data_offset=3;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h2955901066011100A2A8A3AB99518B12A9412A6820120D211ABB0FA388F8F8A4),
    .INIT_01(256'h66002F923C0CC13729201106510C305490A0509AF8A1114E10A22E6332D329A5),
    .INIT_02(256'h99396795B4BF562D15DD5DD643282CA4205744499268260073ABE0EA2A080C23),
    .INIT_03(256'h4921AE9F9718758632775096103CC41C00200354CEFCB8BE14CE48AF21650B44),
    .INIT_04(256'h1E6726628430CD341001428C8A4C5D1C24E2605CFED8C475756F121F7BCBA3B2),
    .INIT_05(256'h08E5202CD07A8F36F1E52BA4696DC04796FD449A6C221AF9004C2B24FD112824),
    .INIT_06(256'h75F06CC44A11872D2B61810F28047025EF296F54B56B37DA81561C1CD6C92700),
    .INIT_07(256'h36FE3E01B8F118F91B1A81854E149A36A60BCC93205C20AC0966C35D944C4FAB),
    .INIT_08(256'hD7FFDCB1A0F06D5849D51168A003568EBBC722FA7EF5D1A90796F12E41F8E020),
    .INIT_09(256'h6EEBAC6590E409EE2F81195E310598B0054E99BB0FA952FA7323E2F0E2B84015),
    .INIT_0A(256'hBDE0918133170B30D82EFDDFEEFCBEBF9BFC7EFCDD70A22E58C4379921BF8388),
    .INIT_0B(256'h9D70F4FC555C2FC3F966045AAAE2949896C1842C0C477435C9E9969D69270EC8),
    .INIT_0C(256'hD166343B88A519149EFDCF23D826223153106CFA934A2B1A1618914F4FF88F84),
    .INIT_0D(256'hFBF661172E3F9F5F44C556E47D9F82FCBF3DDB5BF1DCB78E615CCE588E99CB9D),
    .INIT_0E(256'hC1F759F471BFFFFF19E124FF0FFFF2C63CE79A1B049094E2F99675AD04E72FD7),
    .INIT_0F(256'hD2C02288830A096710E179F77D82026F64A0520A8232A424C0A7840E61EDDB0C),
    .INIT_10(256'hA0001FC40440A4A2F4D0433DB5923622004EBB258C5CEC54D9823307F626537C),
    .INIT_11(256'h776839A304497A936DBB24FBF64968321441CEA996C3000E7126204DFA811488),
    .INIT_12(256'h7E9941BE26FA1F2406264CC5E37A98A81769DB4808666E82426EEC92565DC98B),
    .INIT_13(256'h9CBF4D304384E0B43D4C292DD58C8972FD43A4619CD200CA75602CB92B0A1210),
    .INIT_14(256'hA81456465A1331CD54D94A9E6E51489846131DF0674861E8E5F8FFE3FF5283B4),
    .INIT_15(256'h8F6C603D4B7DF6D95CCA004155B610A2050D10400553605027DFF929C7BE6D79),
    .INIT_16(256'h82288AD4AF18F34600509EB7302225610BC585CAB401014674D3F012AE2B9631),
    .INIT_17(256'hC5C822491EA5F7A5F7F1DEDC7D7F688AC67D6B88D6DA5AA86EEDCF5B06FC8D2A),
    .INIT_18(256'hA5DA1C3EFDA167BE6A8C1816635DF8199E8E361C3A54586406C514040D81410C),
    .INIT_19(256'h8358B1300FECD62885848328C1AD9C99086A262199D19B5B1E70041003020405),
    .INIT_1A(256'hBB3B7214543CC06019C6E11B23C9991731411AD484FB39950B2F0053553C2621),
    .INIT_1B(256'h6FEB68C0F7E0F02082C7E0BFB4FE0FE5F887AAFF17BA1FD7D9B5BCB88C2ACD63),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFF1D801092F6D68B9696884102AA2EC27E98BEF1E56),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_003 (
    .addra(addra),
    .clka(clka),
    .dia({open_n252,open_n253,open_n254,open_n255,open_n256,open_n257,open_n258,1'b0,open_n259}),
    .rsta(rsta),
    .doa({open_n274,open_n275,open_n276,open_n277,open_n278,open_n279,open_n280,open_n281,doa[3]}));
  // address_offset=0;data_offset=4;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h82382A88E04B06401C33236F50554A25C8C19429603A342070C24C2882F8FAA3),
    .INIT_01(256'h89D6D04C80A02248D65D62D1A411C4C82BBBF9EBABFBCA806D0F10842B009427),
    .INIT_02(256'h407FBF8082B7C7D2C8AA0820A04500888B8880A26607D8BC87C21704C462810C),
    .INIT_03(256'hCB20068F741005040044C01602000B1C00205311FAEFAEF904CC94884E922481),
    .INIT_04(256'h3444214029202805B2A64008680A51AB230C9CAA3050D902650B8C0018E81192),
    .INIT_05(256'h54A32D846D44831600CF8AA719EDC4779EBD6C524C8C823203412A2490240940),
    .INIT_06(256'h3645D40C5B64D02B61000F6B2858652C234AD2A4320A9191012000051088B2F8),
    .INIT_07(256'h68402F121020010C1015088004D4000700A2E20027C407B6D3070A880C080411),
    .INIT_08(256'hBC83D800058081D00A0924AC324FC5D8DD01C0440F87C02035A900A54A3A504E),
    .INIT_09(256'h1009642415AC016B06091004D0080104442810FE20500404917D46B50415865C),
    .INIT_0A(256'h04214B4CCF32088741601A410902206400C0294005C70CD1B281A4D0A002A45E),
    .INIT_0B(256'h61ADA502E0CD03169C811A010660E46457864163620D000523460D069762214B),
    .INIT_0C(256'h03D4A76F9208A009E100D40024C8C86DD248A0805068402074CB4BA005032052),
    .INIT_0D(256'h4C9802481802007801AC08508600FC87298843988922843000E044F893BDA230),
    .INIT_0E(256'h660DAB01C24106086306800132521CC320BEB6E6A0EB605BA3BED348355C14A8),
    .INIT_0F(256'h191518DA0455239C55A561844D5A8813C24C80442D24840080146204C3091628),
    .INIT_10(256'h0000409A0000046A4B25100942086987AA6D82DA5C11031F054AA5A811449231),
    .INIT_11(256'h445A222200931D054402DC4839B0692CD08C80ECCA90521184082DB4492D0198),
    .INIT_12(256'h402019079814A004C29019B0E0500185003000D2D044406A5488000599111B4C),
    .INIT_13(256'h306070480E10123A2CCCA13A174D90C11C8D6F9B6200010770991A2D1446EC84),
    .INIT_14(256'hA841704B1786BA7828B29856EEB605F71D4FB22FD2E49A678294A41690C04E60),
    .INIT_15(256'h7A5AC4431A7FA652D1A832611F0D3ADC4493659ED42E456047FB031AA1FE940A),
    .INIT_16(256'h8E1028001000091D288132D2908C2383A6334F40EC643776CFFFF3DDA23C0CE7),
    .INIT_17(256'h722739BF636D0867341B232B4B82D867F33C0B297DE921C0CCCC760E4D96CFA1),
    .INIT_18(256'hD13D339DD104CDC6EE1264CC7B5EFA34C9E6EEE7255335C0DA1827075269BC87),
    .INIT_19(256'hD66346C00F9889C60E936C9BC274E6A6B33806DA367756CEB6840002019CF155),
    .INIT_1A(256'h64241234740CD735F4FD36A4D6624CEA5AB94D8E911C81990BD010165D6CC8CA),
    .INIT_1B(256'hD0E36010A050A20529C72A783048A482968A11243D14115DDF31C691362A6FDA),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFE8194D0005FE7317977040A89D3D0D0241313D57C7),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_004 (
    .addra(addra),
    .clka(clka),
    .dia({open_n313,open_n314,open_n315,open_n316,open_n317,open_n318,open_n319,1'b0,open_n320}),
    .rsta(rsta),
    .doa({open_n335,open_n336,open_n337,open_n338,open_n339,open_n340,open_n341,open_n342,doa[4]}));
  // address_offset=0;data_offset=5;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'hEFFC7F41C1FF402130541DA988270255E8EDB4A0C6425420384026118AFAFA87),
    .INIT_01(256'h000000000000000000000000000000001544005100100143FFFFE3FFFFE0FF7F),
    .INIT_02(256'h001B248A80002A8822822AAA0882111004000000000000000381E00202000000),
    .INIT_03(256'h000C81D39C0C45208855FD1E5E09EF5D00200100630005510466008000030000),
    .INIT_04(256'h97F5FBC63C7E3F8565FB312447080C2B0B0628023013E0A3570B304010CD1404),
    .INIT_05(256'h422301A5426C2A8F80C662E3D463C0418E1C6C561D0E0631593DB91244B367EC),
    .INIT_06(256'h3805D48C5744D0F92900274B18218605294A52A5330891918D2004055080B203),
    .INIT_07(256'h85403C05542BCC1951EA0292A4744A8413C5C549A3060624C71D74890EA08099),
    .INIT_08(256'h90829A40C41662C8468C92BDB947948AA85D3514EF8DF2182D001751EAB9513C),
    .INIT_09(256'h125D642E548EE06201D2D3A0DBC0400173488D13A148A7140616B48E02022005),
    .INIT_0A(256'h842D4B110B300BBC057018EB590A410580C261482509554A908822935DC21C5A),
    .INIT_0B(256'h8D24AC02C9E003123AA14EEB4F018C005E802523FFF4080D0B5B81100562234B),
    .INIT_0C(256'h0A64222B89001819E101CC6E9115518750280089A83D50FFF50E5921AC0D5009),
    .INIT_0D(256'hD9B780A163BA80B8022DE9424480A58C6358C014874908382A00055303B146B4),
    .INIT_0E(256'h93558901D41000806A47940416D20252A98717508B838951A9C4DF7A9D51B4BA),
    .INIT_0F(256'h5E3F109E70F10040558AEB8534E0E6177E42EB2DF8267312434498F15548C849),
    .INIT_10(256'hD77742A8EEDDFC754007910ABA8120A68B0499015CC8CD18217560FF6204C849),
    .INIT_11(256'h53292BB992CB05C85499D04804040DA4D6C0F18AABAAFF281855E4004925803D),
    .INIT_12(256'h5AB489102AD0075F590262000BD45C3F8243EAE1CF5B4475D20A7049B494C978),
    .INIT_13(256'h0421200008045900625D9FC8050CB8103801A0080403BC823B092022C006D006),
    .INIT_14(256'hC84002E77298924C759C1B83324246117189047416C14110209024469010482C),
    .INIT_15(256'hE34001002B24879C663BDD81DC2062100221A00C959867102249700100927D8C),
    .INIT_16(256'h9425535EE9DEEB708C980236B0B00341F860478BAC0DC722649179CA82918E73),
    .INIT_17(256'h6244B56DA0820804602156B840715953A26D8E40905E15066EEE9768B1A2F6AC),
    .INIT_18(256'h85EFA2B1E88F14B332A92DFA0F509A0081D0AB840663E71728E0C20408222844),
    .INIT_19(256'h90C428000FEF9DA00220480E81258C800013BB110D7154880119009442F193FC),
    .INIT_1A(256'h0880056314022209C07008104000039563E9A156552A00C9190831086C851518),
    .INIT_1B(256'hBF408190A850A937FBD63EF0B649F4A092D208A430101F7557B5814E5012CB08),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFE81B050009DAC55EBC11A6FD98182C324255A9150C),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_005 (
    .addra(addra),
    .clka(clka),
    .dia({open_n374,open_n375,open_n376,open_n377,open_n378,open_n379,open_n380,1'b0,open_n381}),
    .rsta(rsta),
    .doa({open_n396,open_n397,open_n398,open_n399,open_n400,open_n401,open_n402,open_n403,doa[5]}));
  // address_offset=0;data_offset=6;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h13FE43BE21EF990C828CADA1810599075940266C4A06959776FBEDBFB1F9F995),
    .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD400004101015501FDBF73F77BF0FFB0),
    .INIT_02(256'hF24B2C8A0802AA0AA20A082A077DEEEFFBFFFFFFFFFFFFFFFC7E1FFDFDFFFFFF),
    .INIT_03(256'h0000135AA80594F658337AD41F0CCF8C249001573503604612EED27FFFFCFFFF),
    .INIT_04(256'hEB73A470ED80CF1220A71761E32404C72E619EE6C6C8C4308967021B73298200),
    .INIT_05(256'h60C5BD3DA1FE65BE36EC65E27CE7D55696C5C89B6C0858C8C019288018200142),
    .INIT_06(256'hBB9D18CA1BD85B9DA46D83276BE41394A7395B34B06303D800B6D8DC86440100),
    .INIT_07(256'h972C8F1DC998C59CC8953900F622039581E3C3C0961ECC2E4970EAEDB56EF300),
    .INIT_08(256'h125DFE106270244322C0004C70E286E88FC0F73630B6DD0935B871A24C586917),
    .INIT_09(256'hCB6ABC0A0834246692DB48B348EC2093516405DBB673B5664E2C3647604E6034),
    .INIT_0A(256'h318072322C234001B65769652DB12D9232DBA4D1B73DF766E6439048A4590DD4),
    .INIT_0B(256'hB0383764AE476C60DE4CC224723719B206D95603EF78BB3262363362B6506D82),
    .INIT_0C(256'hC384A527C06C83312DB2C4E25B3777BDD90436B8D10998FEFB217096B4B5CB38),
    .INIT_0D(256'h6AD74A25E78936DBC6C8672E1D365295A52B48F7B12C91A315DF52B2862DA256),
    .INIT_0E(256'h706D90711ADB76DB5374C1D9DB5971684C08BBDBF4BA183C86D485AC5777F66D),
    .INIT_0F(256'h6E75589207530427D91524B31068A0DBBF7EB803AD90317A0772390649244304),
    .INIT_10(256'h71116C6E220474AB265DE667593D32D44A36886D904450EA6CEB3BA93112036F),
    .INIT_11(256'h31051AA880A227832508C26B46D89D168083D6B332B1D3077BB330DB24C03268),
    .INIT_12(256'h252C2C8BEE0B09A77A6E2EEC88CDC6DDB1B1357FFF3F23AA582620C136CC6C89),
    .INIT_13(256'hC9B6259241F9FC8DA32FDD24F9C233265A47936DDDE34E62DE6F0595098AA715),
    .INIT_14(256'hA98A9CD61983776903BF6D9AAB1908D9039DDDC6615E6D8A4EC93D8ACB2681B0),
    .INIT_15(256'h0E67603FE6B6C185E2C8C4604593A036034C36FC841115201B6D949CA6DB546A),
    .INIT_16(256'hC40AA8C62FC63B1240C00D1103072D64D1A5D720B498494556D31ED12FAED4A5),
    .INIT_17(256'hA7DED76D92316DBDA5DC8A6C98D628CB8F0C52C8D21C5EFF55550E1982C8C222),
    .INIT_18(256'hD00C46D6CC57664AAA2FB0010C22921B335BBB1C8CE40C3104645D05E59E59F7),
    .INIT_19(256'h735CBC300F999B91C34DF962D5B41019DEC88B3DEDFC9999D87A009002E29752),
    .INIT_1A(256'hBBCB5311242B4ED38B22D3DB7B49B5D5AEAD116C88FB6891122D11534D17773F),
    .INIT_1B(256'hA00848EA286A2C8D28C6EA363167B64ECBBB99B3124E13B793756A629E0A192C),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFEDC56025926B4DFCE25891A8A2928C0B24DFCD4694),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_006 (
    .addra(addra),
    .clka(clka),
    .dia({open_n435,open_n436,open_n437,open_n438,open_n439,open_n440,open_n441,1'b0,open_n442}),
    .rsta(rsta),
    .doa({open_n457,open_n458,open_n459,open_n460,open_n461,open_n462,open_n463,open_n464,doa[6]}));
  // address_offset=0;data_offset=7;depth=8192;width=1;num_section=1;width_per_section=1;section_size=8;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000001B04E68DAA51B1CD9BC2839A6664100F04B3F3EFFCFD99F9F99D),
    .INIT_01(256'h1084810908222445224108148912111240104301540524400000000000000000),
    .INIT_02(256'h0002400A0BE8082A2AA0AA88B1042222489088924924924927A7E24454484211),
    .INIT_03(256'h001A131E682591F6D87788700000002F2490015A9ECEAE8C1088D2C000000000),
    .INIT_04(256'hE806050CC5B061170C059771F06C25EF6F339C66424ECD3D8A2F66996309E200),
    .INIT_05(256'h60E61735A1BCEEB4178E6F4745AD1516B4E5B8DA6B1BD8CCE4876EC90E68D03A),
    .INIT_06(256'hA9BF1CD99BDF59B6CC65906229EF33B4A5295B35AD61E29E98B6585886471D06),
    .INIT_07(256'hB764989DDDBEE59DDC813B08F707B1B4EDF9DBF6931A46024A70E0E49826F3E6),
    .INIT_08(256'h16CCD7837A7D24A12AF648D774FA86E88FE1C733B096982835F83D070E542D97),
    .INIT_09(256'hDB6BC00A0E39A4EE921B5EB36EEC6093DD6C25A5B2739D264E0C06D7204A631E),
    .INIT_0A(256'hB1987E776EE3344097D729673D9165B6B799A4859C3DF766E2E1BC5E064B4DF6),
    .INIT_0B(256'h90363427AE8F2C38D6CDE72C7473399784CB178000019930363E332297CC6FB6),
    .INIT_0C(256'h6364A70D642C833F2C92A49ADF3773BCDB8C339C8120D80003633CB29495D938),
    .INIT_0D(256'hEAF402ADE7CB36D186FA6F6F1936F7BCAF69C856916D90EB901956C24D65F066),
    .INIT_0E(256'h1929B42B1ADB26D9CB6DD1C9C81B63FCC48BAD5BE03E9A7D070186724377F6FD),
    .INIT_0F(256'h6EF05831060304365F304D379269B0CA3F7BBC5384B1097B0736B9028A2E638E),
    .INIT_10(256'h799964EF332640C16E48966E1B3D326CE6094E6CF066508AEDE1018128162369),
    .INIT_11(256'h79853EEE89AB27A3644ED66B46C8973789A1529998A1818F691710C96DB2B273),
    .INIT_12(256'h606E0DC0EF1B08033A6F2EE49C9CE6C0B80021BFF37C70E0382F2061A65E6CC1),
    .INIT_13(256'hC9B22697F1B9ED85A36B100CD64A3326DA469B65D8800EE06B66849009AD975D),
    .INIT_14(256'h11AA9B878B63868197A0721444D908DB931DDDC3799E658A4EDB388CD92731BF),
    .INIT_15(256'h066F62386C0019A582E4D5026097843233043676A21BA9941000A480A524A251),
    .INIT_16(256'hC04804E12FE73696D0209D99C3422E65F385B29C189A4E8800030EE135C1A108),
    .INIT_17(256'hAFDED76EB1B12CB5A4819AED99D630D9459A54C8C38A5F0F99998D93A7600012),
    .INIT_18(256'hD00C06D68CD366C4442FB0030C06B6191359B9950EE404794EED59A0EDBE5BE9),
    .INIT_19(256'h731DBD38C3634043434CFB225C9E391BCECCC93CE5ADDCB3D87A0010E272A602),
    .INIT_1A(256'hBBDB9D8CB04B4E53D96651CB7B51944E440E303922232625146CC1E38637377F),
    .INIT_1B(256'h900848CA280A28C88084C026296F16CED91BEEB7C2CF0C6A28684A62190F196D),
    .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFEDCF382492694CCC52C899182292884B64CCCD4694),
    .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x8_sub_000000_007 (
    .addra(addra),
    .clka(clka),
    .dia({open_n496,open_n497,open_n498,open_n499,open_n500,open_n501,open_n502,1'b0,open_n503}),
    .rsta(rsta),
    .doa({open_n518,open_n519,open_n520,open_n521,open_n522,open_n523,open_n524,open_n525,doa[7]}));

endmodule 

