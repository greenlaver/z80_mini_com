//
// Microsoft-BASIC ROM for Z80
//
module basic_microm(n_rst, clk, ce, oe, addr, data);

input        n_rst, clk;
input        ce, oe;
input  [12:0] addr;
output [7:0] data;

reg [7:0] data_buf;

always @(posedge clk or negedge n_rst) begin
	if(!n_rst) begin
		data_buf <= 8'hzz;
	end
	else begin
		case (addr)
			13'h0000: data_buf = 8'hf3;
			13'h0001: data_buf = 8'h31;
			13'h0002: data_buf = 8'hed;
			13'h0003: data_buf = 8'h80;
			13'h0004: data_buf = 8'hc3;
			13'h0005: data_buf = 8'h1b;
			13'h0006: data_buf = 8'h00;
			13'h0007: data_buf = 8'hff;
			13'h0008: data_buf = 8'hc3;
			13'h0009: data_buf = 8'h36;
			13'h000a: data_buf = 8'h00;
			13'h000b: data_buf = 8'hff;
			13'h000c: data_buf = 8'hff;
			13'h000d: data_buf = 8'hff;
			13'h000e: data_buf = 8'hff;
			13'h000f: data_buf = 8'hff;
			13'h0010: data_buf = 8'hc3;
			13'h0011: data_buf = 8'h22;
			13'h0012: data_buf = 8'h00;
			13'h0013: data_buf = 8'hff;
			13'h0014: data_buf = 8'hff;
			13'h0015: data_buf = 8'hff;
			13'h0016: data_buf = 8'hff;
			13'h0017: data_buf = 8'hff;
			13'h0018: data_buf = 8'hc3;
			13'h0019: data_buf = 8'h31;
			13'h001a: data_buf = 8'h00;
			13'h001b: data_buf = 8'haf;
			13'h001c: data_buf = 8'hc3;
			13'h001d: data_buf = 8'h41;
			13'h001e: data_buf = 8'h00;
			13'h001f: data_buf = 8'hfb;
			13'h0020: data_buf = 8'hed;
			13'h0021: data_buf = 8'h4d;
			13'h0022: data_buf = 8'hc5;
			13'h0023: data_buf = 8'hd5;
			13'h0024: data_buf = 8'he5;
			13'h0025: data_buf = 8'hdb;
			13'h0026: data_buf = 8'h85;
			13'h0027: data_buf = 8'hcb;
			13'h0028: data_buf = 8'h4f;
			13'h0029: data_buf = 8'h28;
			13'h002a: data_buf = 8'hfa;
			13'h002b: data_buf = 8'hdb;
			13'h002c: data_buf = 8'h84;
			13'h002d: data_buf = 8'he1;
			13'h002e: data_buf = 8'hd1;
			13'h002f: data_buf = 8'hc1;
			13'h0030: data_buf = 8'hc9;
			13'h0031: data_buf = 8'hdb;
			13'h0032: data_buf = 8'h85;
			13'h0033: data_buf = 8'hcb;
			13'h0034: data_buf = 8'h4f;
			13'h0035: data_buf = 8'hc9;
			13'h0036: data_buf = 8'hf5;
			13'h0037: data_buf = 8'hdb;
			13'h0038: data_buf = 8'h85;
			13'h0039: data_buf = 8'hcb;
			13'h003a: data_buf = 8'h47;
			13'h003b: data_buf = 8'h28;
			13'h003c: data_buf = 8'hfa;
			13'h003d: data_buf = 8'hf1;
			13'h003e: data_buf = 8'hd3;
			13'h003f: data_buf = 8'h84;
			13'h0040: data_buf = 8'hc9;
			13'h0041: data_buf = 8'hc3;
			13'h0042: data_buf = 8'h47;
			13'h0043: data_buf = 8'h00;
			13'h0044: data_buf = 8'hc3;
			13'h0045: data_buf = 8'hbc;
			13'h0046: data_buf = 8'h00;
			13'h0047: data_buf = 8'hc3;
			13'h0048: data_buf = 8'h4e;
			13'h0049: data_buf = 8'h00;
			13'h004a: data_buf = 8'hff;
			13'h004b: data_buf = 8'h08;
			13'h004c: data_buf = 8'h75;
			13'h004d: data_buf = 8'h10;
			13'h004e: data_buf = 8'h21;
			13'h004f: data_buf = 8'h45;
			13'h0050: data_buf = 8'h80;
			13'h0051: data_buf = 8'hf9;
			13'h0052: data_buf = 8'hc3;
			13'h0053: data_buf = 8'h90;
			13'h0054: data_buf = 8'h1c;
			13'h0055: data_buf = 8'h11;
			13'h0056: data_buf = 8'h26;
			13'h0057: data_buf = 8'h03;
			13'h0058: data_buf = 8'h06;
			13'h0059: data_buf = 8'h63;
			13'h005a: data_buf = 8'h21;
			13'h005b: data_buf = 8'h45;
			13'h005c: data_buf = 8'h80;
			13'h005d: data_buf = 8'h1a;
			13'h005e: data_buf = 8'h77;
			13'h005f: data_buf = 8'h23;
			13'h0060: data_buf = 8'h13;
			13'h0061: data_buf = 8'h05;
			13'h0062: data_buf = 8'hc2;
			13'h0063: data_buf = 8'h5d;
			13'h0064: data_buf = 8'h00;
			13'h0065: data_buf = 8'hf9;
			13'h0066: data_buf = 8'hcd;
			13'h0067: data_buf = 8'h27;
			13'h0068: data_buf = 8'h05;
			13'h0069: data_buf = 8'hcd;
			13'h006a: data_buf = 8'hf5;
			13'h006b: data_buf = 8'h0a;
			13'h006c: data_buf = 8'h32;
			13'h006d: data_buf = 8'hef;
			13'h006e: data_buf = 8'h80;
			13'h006f: data_buf = 8'h32;
			13'h0070: data_buf = 8'h3e;
			13'h0071: data_buf = 8'h81;
			13'h0072: data_buf = 8'h21;
			13'h0073: data_buf = 8'ha2;
			13'h0074: data_buf = 8'h81;
			13'h0075: data_buf = 8'h23;
			13'h0076: data_buf = 8'h7c;
			13'h0077: data_buf = 8'hb5;
			13'h0078: data_buf = 8'hca;
			13'h0079: data_buf = 8'h84;
			13'h007a: data_buf = 8'h00;
			13'h007b: data_buf = 8'h7e;
			13'h007c: data_buf = 8'h47;
			13'h007d: data_buf = 8'h2f;
			13'h007e: data_buf = 8'h77;
			13'h007f: data_buf = 8'hbe;
			13'h0080: data_buf = 8'h70;
			13'h0081: data_buf = 8'hca;
			13'h0082: data_buf = 8'h75;
			13'h0083: data_buf = 8'h00;
			13'h0084: data_buf = 8'h2b;
			13'h0085: data_buf = 8'h11;
			13'h0086: data_buf = 8'ha1;
			13'h0087: data_buf = 8'h81;
			13'h0088: data_buf = 8'hcd;
			13'h0089: data_buf = 8'hbd;
			13'h008a: data_buf = 8'h06;
			13'h008b: data_buf = 8'hda;
			13'h008c: data_buf = 8'hc5;
			13'h008d: data_buf = 8'h00;
			13'h008e: data_buf = 8'h11;
			13'h008f: data_buf = 8'hce;
			13'h0090: data_buf = 8'hff;
			13'h0091: data_buf = 8'h22;
			13'h0092: data_buf = 8'hf4;
			13'h0093: data_buf = 8'h80;
			13'h0094: data_buf = 8'h19;
			13'h0095: data_buf = 8'h22;
			13'h0096: data_buf = 8'h9f;
			13'h0097: data_buf = 8'h80;
			13'h0098: data_buf = 8'hcd;
			13'h0099: data_buf = 8'h02;
			13'h009a: data_buf = 8'h05;
			13'h009b: data_buf = 8'h2a;
			13'h009c: data_buf = 8'h9f;
			13'h009d: data_buf = 8'h80;
			13'h009e: data_buf = 8'h11;
			13'h009f: data_buf = 8'hef;
			13'h00a0: data_buf = 8'hff;
			13'h00a1: data_buf = 8'h19;
			13'h00a2: data_buf = 8'h11;
			13'h00a3: data_buf = 8'h3e;
			13'h00a4: data_buf = 8'h81;
			13'h00a5: data_buf = 8'h7d;
			13'h00a6: data_buf = 8'h93;
			13'h00a7: data_buf = 8'h6f;
			13'h00a8: data_buf = 8'h7c;
			13'h00a9: data_buf = 8'h9a;
			13'h00aa: data_buf = 8'h67;
			13'h00ab: data_buf = 8'he5;
			13'h00ac: data_buf = 8'h21;
			13'h00ad: data_buf = 8'hdd;
			13'h00ae: data_buf = 8'h00;
			13'h00af: data_buf = 8'hcd;
			13'h00b0: data_buf = 8'h93;
			13'h00b1: data_buf = 8'h11;
			13'h00b2: data_buf = 8'he1;
			13'h00b3: data_buf = 8'hcd;
			13'h00b4: data_buf = 8'h36;
			13'h00b5: data_buf = 8'h18;
			13'h00b6: data_buf = 8'h21;
			13'h00b7: data_buf = 8'hce;
			13'h00b8: data_buf = 8'h00;
			13'h00b9: data_buf = 8'hcd;
			13'h00ba: data_buf = 8'h93;
			13'h00bb: data_buf = 8'h11;
			13'h00bc: data_buf = 8'h31;
			13'h00bd: data_buf = 8'hab;
			13'h00be: data_buf = 8'h80;
			13'h00bf: data_buf = 8'hcd;
			13'h00c0: data_buf = 8'h27;
			13'h00c1: data_buf = 8'h05;
			13'h00c2: data_buf = 8'hc3;
			13'h00c3: data_buf = 8'h40;
			13'h00c4: data_buf = 8'h04;
			13'h00c5: data_buf = 8'h21;
			13'h00c6: data_buf = 8'h14;
			13'h00c7: data_buf = 8'h01;
			13'h00c8: data_buf = 8'hcd;
			13'h00c9: data_buf = 8'h93;
			13'h00ca: data_buf = 8'h11;
			13'h00cb: data_buf = 8'hc3;
			13'h00cc: data_buf = 8'hcb;
			13'h00cd: data_buf = 8'h00;
			13'h00ce: data_buf = 8'h20;
			13'h00cf: data_buf = 8'h42;
			13'h00d0: data_buf = 8'h79;
			13'h00d1: data_buf = 8'h74;
			13'h00d2: data_buf = 8'h65;
			13'h00d3: data_buf = 8'h73;
			13'h00d4: data_buf = 8'h20;
			13'h00d5: data_buf = 8'h66;
			13'h00d6: data_buf = 8'h72;
			13'h00d7: data_buf = 8'h65;
			13'h00d8: data_buf = 8'h65;
			13'h00d9: data_buf = 8'h0d;
			13'h00da: data_buf = 8'h0a;
			13'h00db: data_buf = 8'h00;
			13'h00dc: data_buf = 8'h00;
			13'h00dd: data_buf = 8'h5a;
			13'h00de: data_buf = 8'h38;
			13'h00df: data_buf = 8'h30;
			13'h00e0: data_buf = 8'h20;
			13'h00e1: data_buf = 8'h42;
			13'h00e2: data_buf = 8'h41;
			13'h00e3: data_buf = 8'h53;
			13'h00e4: data_buf = 8'h49;
			13'h00e5: data_buf = 8'h43;
			13'h00e6: data_buf = 8'h20;
			13'h00e7: data_buf = 8'h56;
			13'h00e8: data_buf = 8'h65;
			13'h00e9: data_buf = 8'h72;
			13'h00ea: data_buf = 8'h20;
			13'h00eb: data_buf = 8'h34;
			13'h00ec: data_buf = 8'h2e;
			13'h00ed: data_buf = 8'h37;
			13'h00ee: data_buf = 8'h62;
			13'h00ef: data_buf = 8'h0d;
			13'h00f0: data_buf = 8'h0a;
			13'h00f1: data_buf = 8'h43;
			13'h00f2: data_buf = 8'h6f;
			13'h00f3: data_buf = 8'h70;
			13'h00f4: data_buf = 8'h79;
			13'h00f5: data_buf = 8'h72;
			13'h00f6: data_buf = 8'h69;
			13'h00f7: data_buf = 8'h67;
			13'h00f8: data_buf = 8'h68;
			13'h00f9: data_buf = 8'h74;
			13'h00fa: data_buf = 8'h20;
			13'h00fb: data_buf = 8'h28;
			13'h00fc: data_buf = 8'h43;
			13'h00fd: data_buf = 8'h29;
			13'h00fe: data_buf = 8'h20;
			13'h00ff: data_buf = 8'h31;
			13'h0100: data_buf = 8'h39;
			13'h0101: data_buf = 8'h37;
			13'h0102: data_buf = 8'h38;
			13'h0103: data_buf = 8'h20;
			13'h0104: data_buf = 8'h62;
			13'h0105: data_buf = 8'h79;
			13'h0106: data_buf = 8'h20;
			13'h0107: data_buf = 8'h4d;
			13'h0108: data_buf = 8'h69;
			13'h0109: data_buf = 8'h63;
			13'h010a: data_buf = 8'h72;
			13'h010b: data_buf = 8'h6f;
			13'h010c: data_buf = 8'h73;
			13'h010d: data_buf = 8'h6f;
			13'h010e: data_buf = 8'h66;
			13'h010f: data_buf = 8'h74;
			13'h0110: data_buf = 8'h0d;
			13'h0111: data_buf = 8'h0a;
			13'h0112: data_buf = 8'h00;
			13'h0113: data_buf = 8'h00;
			13'h0114: data_buf = 8'h4d;
			13'h0115: data_buf = 8'h65;
			13'h0116: data_buf = 8'h6d;
			13'h0117: data_buf = 8'h6f;
			13'h0118: data_buf = 8'h72;
			13'h0119: data_buf = 8'h79;
			13'h011a: data_buf = 8'h20;
			13'h011b: data_buf = 8'h73;
			13'h011c: data_buf = 8'h69;
			13'h011d: data_buf = 8'h7a;
			13'h011e: data_buf = 8'h65;
			13'h011f: data_buf = 8'h20;
			13'h0120: data_buf = 8'h6e;
			13'h0121: data_buf = 8'h6f;
			13'h0122: data_buf = 8'h74;
			13'h0123: data_buf = 8'h20;
			13'h0124: data_buf = 8'h65;
			13'h0125: data_buf = 8'h6e;
			13'h0126: data_buf = 8'h6f;
			13'h0127: data_buf = 8'h75;
			13'h0128: data_buf = 8'h67;
			13'h0129: data_buf = 8'h68;
			13'h012a: data_buf = 8'h0d;
			13'h012b: data_buf = 8'h0a;
			13'h012c: data_buf = 8'h54;
			13'h012d: data_buf = 8'h68;
			13'h012e: data_buf = 8'h65;
			13'h012f: data_buf = 8'h20;
			13'h0130: data_buf = 8'h73;
			13'h0131: data_buf = 8'h79;
			13'h0132: data_buf = 8'h73;
			13'h0133: data_buf = 8'h74;
			13'h0134: data_buf = 8'h65;
			13'h0135: data_buf = 8'h6d;
			13'h0136: data_buf = 8'h20;
			13'h0137: data_buf = 8'h69;
			13'h0138: data_buf = 8'h73;
			13'h0139: data_buf = 8'h20;
			13'h013a: data_buf = 8'h73;
			13'h013b: data_buf = 8'h74;
			13'h013c: data_buf = 8'h6f;
			13'h013d: data_buf = 8'h70;
			13'h013e: data_buf = 8'h70;
			13'h013f: data_buf = 8'h65;
			13'h0140: data_buf = 8'h64;
			13'h0141: data_buf = 8'h2e;
			13'h0142: data_buf = 8'h0d;
			13'h0143: data_buf = 8'h0a;
			13'h0144: data_buf = 8'h00;
			13'h0145: data_buf = 8'h00;
			13'h0146: data_buf = 8'hab;
			13'h0147: data_buf = 8'h16;
			13'h0148: data_buf = 8'h6f;
			13'h0149: data_buf = 8'h17;
			13'h014a: data_buf = 8'hc1;
			13'h014b: data_buf = 8'h16;
			13'h014c: data_buf = 8'h48;
			13'h014d: data_buf = 8'h80;
			13'h014e: data_buf = 8'h53;
			13'h014f: data_buf = 8'h10;
			13'h0150: data_buf = 8'hd8;
			13'h0151: data_buf = 8'h13;
			13'h0152: data_buf = 8'h81;
			13'h0153: data_buf = 8'h10;
			13'h0154: data_buf = 8'h35;
			13'h0155: data_buf = 8'h19;
			13'h0156: data_buf = 8'h14;
			13'h0157: data_buf = 8'h1a;
			13'h0158: data_buf = 8'h50;
			13'h0159: data_buf = 8'h15;
			13'h015a: data_buf = 8'h83;
			13'h015b: data_buf = 8'h19;
			13'h015c: data_buf = 8'h89;
			13'h015d: data_buf = 8'h1a;
			13'h015e: data_buf = 8'h8f;
			13'h015f: data_buf = 8'h1a;
			13'h0160: data_buf = 8'hf0;
			13'h0161: data_buf = 8'h1a;
			13'h0162: data_buf = 8'h05;
			13'h0163: data_buf = 8'h1b;
			13'h0164: data_buf = 8'h2c;
			13'h0165: data_buf = 8'h14;
			13'h0166: data_buf = 8'h70;
			13'h0167: data_buf = 8'h1b;
			13'h0168: data_buf = 8'h96;
			13'h0169: data_buf = 8'h80;
			13'h016a: data_buf = 8'h05;
			13'h016b: data_buf = 8'h13;
			13'h016c: data_buf = 8'h1d;
			13'h016d: data_buf = 8'h11;
			13'h016e: data_buf = 8'h9f;
			13'h016f: data_buf = 8'h13;
			13'h0170: data_buf = 8'h14;
			13'h0171: data_buf = 8'h13;
			13'h0172: data_buf = 8'h25;
			13'h0173: data_buf = 8'h13;
			13'h0174: data_buf = 8'h92;
			13'h0175: data_buf = 8'h1b;
			13'h0176: data_buf = 8'h25;
			13'h0177: data_buf = 8'h1c;
			13'h0178: data_buf = 8'h35;
			13'h0179: data_buf = 8'h13;
			13'h017a: data_buf = 8'h65;
			13'h017b: data_buf = 8'h13;
			13'h017c: data_buf = 8'h6f;
			13'h017d: data_buf = 8'h13;
			13'h017e: data_buf = 8'hc5;
			13'h017f: data_buf = 8'h4e;
			13'h0180: data_buf = 8'h44;
			13'h0181: data_buf = 8'hc6;
			13'h0182: data_buf = 8'h4f;
			13'h0183: data_buf = 8'h52;
			13'h0184: data_buf = 8'hce;
			13'h0185: data_buf = 8'h45;
			13'h0186: data_buf = 8'h58;
			13'h0187: data_buf = 8'h54;
			13'h0188: data_buf = 8'hc4;
			13'h0189: data_buf = 8'h41;
			13'h018a: data_buf = 8'h54;
			13'h018b: data_buf = 8'h41;
			13'h018c: data_buf = 8'hc9;
			13'h018d: data_buf = 8'h4e;
			13'h018e: data_buf = 8'h50;
			13'h018f: data_buf = 8'h55;
			13'h0190: data_buf = 8'h54;
			13'h0191: data_buf = 8'hc4;
			13'h0192: data_buf = 8'h49;
			13'h0193: data_buf = 8'h4d;
			13'h0194: data_buf = 8'hd2;
			13'h0195: data_buf = 8'h45;
			13'h0196: data_buf = 8'h41;
			13'h0197: data_buf = 8'h44;
			13'h0198: data_buf = 8'hcc;
			13'h0199: data_buf = 8'h45;
			13'h019a: data_buf = 8'h54;
			13'h019b: data_buf = 8'hc7;
			13'h019c: data_buf = 8'h4f;
			13'h019d: data_buf = 8'h54;
			13'h019e: data_buf = 8'h4f;
			13'h019f: data_buf = 8'hd2;
			13'h01a0: data_buf = 8'h55;
			13'h01a1: data_buf = 8'h4e;
			13'h01a2: data_buf = 8'hc9;
			13'h01a3: data_buf = 8'h46;
			13'h01a4: data_buf = 8'hd2;
			13'h01a5: data_buf = 8'h45;
			13'h01a6: data_buf = 8'h53;
			13'h01a7: data_buf = 8'h54;
			13'h01a8: data_buf = 8'h4f;
			13'h01a9: data_buf = 8'h52;
			13'h01aa: data_buf = 8'h45;
			13'h01ab: data_buf = 8'hc7;
			13'h01ac: data_buf = 8'h4f;
			13'h01ad: data_buf = 8'h53;
			13'h01ae: data_buf = 8'h55;
			13'h01af: data_buf = 8'h42;
			13'h01b0: data_buf = 8'hd2;
			13'h01b1: data_buf = 8'h45;
			13'h01b2: data_buf = 8'h54;
			13'h01b3: data_buf = 8'h55;
			13'h01b4: data_buf = 8'h52;
			13'h01b5: data_buf = 8'h4e;
			13'h01b6: data_buf = 8'hd2;
			13'h01b7: data_buf = 8'h45;
			13'h01b8: data_buf = 8'h4d;
			13'h01b9: data_buf = 8'hd3;
			13'h01ba: data_buf = 8'h54;
			13'h01bb: data_buf = 8'h4f;
			13'h01bc: data_buf = 8'h50;
			13'h01bd: data_buf = 8'hcf;
			13'h01be: data_buf = 8'h55;
			13'h01bf: data_buf = 8'h54;
			13'h01c0: data_buf = 8'hcf;
			13'h01c1: data_buf = 8'h4e;
			13'h01c2: data_buf = 8'hce;
			13'h01c3: data_buf = 8'h55;
			13'h01c4: data_buf = 8'h4c;
			13'h01c5: data_buf = 8'h4c;
			13'h01c6: data_buf = 8'hd7;
			13'h01c7: data_buf = 8'h41;
			13'h01c8: data_buf = 8'h49;
			13'h01c9: data_buf = 8'h54;
			13'h01ca: data_buf = 8'hc4;
			13'h01cb: data_buf = 8'h45;
			13'h01cc: data_buf = 8'h46;
			13'h01cd: data_buf = 8'hd0;
			13'h01ce: data_buf = 8'h4f;
			13'h01cf: data_buf = 8'h4b;
			13'h01d0: data_buf = 8'h45;
			13'h01d1: data_buf = 8'hc4;
			13'h01d2: data_buf = 8'h4f;
			13'h01d3: data_buf = 8'h4b;
			13'h01d4: data_buf = 8'h45;
			13'h01d5: data_buf = 8'hd3;
			13'h01d6: data_buf = 8'h43;
			13'h01d7: data_buf = 8'h52;
			13'h01d8: data_buf = 8'h45;
			13'h01d9: data_buf = 8'h45;
			13'h01da: data_buf = 8'h4e;
			13'h01db: data_buf = 8'hcc;
			13'h01dc: data_buf = 8'h49;
			13'h01dd: data_buf = 8'h4e;
			13'h01de: data_buf = 8'h45;
			13'h01df: data_buf = 8'h53;
			13'h01e0: data_buf = 8'hc3;
			13'h01e1: data_buf = 8'h4c;
			13'h01e2: data_buf = 8'h53;
			13'h01e3: data_buf = 8'hd7;
			13'h01e4: data_buf = 8'h49;
			13'h01e5: data_buf = 8'h44;
			13'h01e6: data_buf = 8'h54;
			13'h01e7: data_buf = 8'h48;
			13'h01e8: data_buf = 8'hcd;
			13'h01e9: data_buf = 8'h4f;
			13'h01ea: data_buf = 8'h4e;
			13'h01eb: data_buf = 8'h49;
			13'h01ec: data_buf = 8'h54;
			13'h01ed: data_buf = 8'h4f;
			13'h01ee: data_buf = 8'h52;
			13'h01ef: data_buf = 8'hd3;
			13'h01f0: data_buf = 8'h45;
			13'h01f1: data_buf = 8'h54;
			13'h01f2: data_buf = 8'hd2;
			13'h01f3: data_buf = 8'h45;
			13'h01f4: data_buf = 8'h53;
			13'h01f5: data_buf = 8'h45;
			13'h01f6: data_buf = 8'h54;
			13'h01f7: data_buf = 8'hd0;
			13'h01f8: data_buf = 8'h52;
			13'h01f9: data_buf = 8'h49;
			13'h01fa: data_buf = 8'h4e;
			13'h01fb: data_buf = 8'h54;
			13'h01fc: data_buf = 8'hc3;
			13'h01fd: data_buf = 8'h4f;
			13'h01fe: data_buf = 8'h4e;
			13'h01ff: data_buf = 8'h54;
			13'h0200: data_buf = 8'hcc;
			13'h0201: data_buf = 8'h49;
			13'h0202: data_buf = 8'h53;
			13'h0203: data_buf = 8'h54;
			13'h0204: data_buf = 8'hc3;
			13'h0205: data_buf = 8'h4c;
			13'h0206: data_buf = 8'h45;
			13'h0207: data_buf = 8'h41;
			13'h0208: data_buf = 8'h52;
			13'h0209: data_buf = 8'hc3;
			13'h020a: data_buf = 8'h4c;
			13'h020b: data_buf = 8'h4f;
			13'h020c: data_buf = 8'h41;
			13'h020d: data_buf = 8'h44;
			13'h020e: data_buf = 8'hc3;
			13'h020f: data_buf = 8'h53;
			13'h0210: data_buf = 8'h41;
			13'h0211: data_buf = 8'h56;
			13'h0212: data_buf = 8'h45;
			13'h0213: data_buf = 8'hce;
			13'h0214: data_buf = 8'h45;
			13'h0215: data_buf = 8'h57;
			13'h0216: data_buf = 8'hd4;
			13'h0217: data_buf = 8'h41;
			13'h0218: data_buf = 8'h42;
			13'h0219: data_buf = 8'h28;
			13'h021a: data_buf = 8'hd4;
			13'h021b: data_buf = 8'h4f;
			13'h021c: data_buf = 8'hc6;
			13'h021d: data_buf = 8'h4e;
			13'h021e: data_buf = 8'hd3;
			13'h021f: data_buf = 8'h50;
			13'h0220: data_buf = 8'h43;
			13'h0221: data_buf = 8'h28;
			13'h0222: data_buf = 8'hd4;
			13'h0223: data_buf = 8'h48;
			13'h0224: data_buf = 8'h45;
			13'h0225: data_buf = 8'h4e;
			13'h0226: data_buf = 8'hce;
			13'h0227: data_buf = 8'h4f;
			13'h0228: data_buf = 8'h54;
			13'h0229: data_buf = 8'hd3;
			13'h022a: data_buf = 8'h54;
			13'h022b: data_buf = 8'h45;
			13'h022c: data_buf = 8'h50;
			13'h022d: data_buf = 8'hab;
			13'h022e: data_buf = 8'had;
			13'h022f: data_buf = 8'haa;
			13'h0230: data_buf = 8'haf;
			13'h0231: data_buf = 8'hde;
			13'h0232: data_buf = 8'hc1;
			13'h0233: data_buf = 8'h4e;
			13'h0234: data_buf = 8'h44;
			13'h0235: data_buf = 8'hcf;
			13'h0236: data_buf = 8'h52;
			13'h0237: data_buf = 8'hbe;
			13'h0238: data_buf = 8'hbd;
			13'h0239: data_buf = 8'hbc;
			13'h023a: data_buf = 8'hd3;
			13'h023b: data_buf = 8'h47;
			13'h023c: data_buf = 8'h4e;
			13'h023d: data_buf = 8'hc9;
			13'h023e: data_buf = 8'h4e;
			13'h023f: data_buf = 8'h54;
			13'h0240: data_buf = 8'hc1;
			13'h0241: data_buf = 8'h42;
			13'h0242: data_buf = 8'h53;
			13'h0243: data_buf = 8'hd5;
			13'h0244: data_buf = 8'h53;
			13'h0245: data_buf = 8'h52;
			13'h0246: data_buf = 8'hc6;
			13'h0247: data_buf = 8'h52;
			13'h0248: data_buf = 8'h45;
			13'h0249: data_buf = 8'hc9;
			13'h024a: data_buf = 8'h4e;
			13'h024b: data_buf = 8'h50;
			13'h024c: data_buf = 8'hd0;
			13'h024d: data_buf = 8'h4f;
			13'h024e: data_buf = 8'h53;
			13'h024f: data_buf = 8'hd3;
			13'h0250: data_buf = 8'h51;
			13'h0251: data_buf = 8'h52;
			13'h0252: data_buf = 8'hd2;
			13'h0253: data_buf = 8'h4e;
			13'h0254: data_buf = 8'h44;
			13'h0255: data_buf = 8'hcc;
			13'h0256: data_buf = 8'h4f;
			13'h0257: data_buf = 8'h47;
			13'h0258: data_buf = 8'hc5;
			13'h0259: data_buf = 8'h58;
			13'h025a: data_buf = 8'h50;
			13'h025b: data_buf = 8'hc3;
			13'h025c: data_buf = 8'h4f;
			13'h025d: data_buf = 8'h53;
			13'h025e: data_buf = 8'hd3;
			13'h025f: data_buf = 8'h49;
			13'h0260: data_buf = 8'h4e;
			13'h0261: data_buf = 8'hd4;
			13'h0262: data_buf = 8'h41;
			13'h0263: data_buf = 8'h4e;
			13'h0264: data_buf = 8'hc1;
			13'h0265: data_buf = 8'h54;
			13'h0266: data_buf = 8'h4e;
			13'h0267: data_buf = 8'hd0;
			13'h0268: data_buf = 8'h45;
			13'h0269: data_buf = 8'h45;
			13'h026a: data_buf = 8'h4b;
			13'h026b: data_buf = 8'hc4;
			13'h026c: data_buf = 8'h45;
			13'h026d: data_buf = 8'h45;
			13'h026e: data_buf = 8'h4b;
			13'h026f: data_buf = 8'hd0;
			13'h0270: data_buf = 8'h4f;
			13'h0271: data_buf = 8'h49;
			13'h0272: data_buf = 8'h4e;
			13'h0273: data_buf = 8'h54;
			13'h0274: data_buf = 8'hcc;
			13'h0275: data_buf = 8'h45;
			13'h0276: data_buf = 8'h4e;
			13'h0277: data_buf = 8'hd3;
			13'h0278: data_buf = 8'h54;
			13'h0279: data_buf = 8'h52;
			13'h027a: data_buf = 8'h24;
			13'h027b: data_buf = 8'hd6;
			13'h027c: data_buf = 8'h41;
			13'h027d: data_buf = 8'h4c;
			13'h027e: data_buf = 8'hc1;
			13'h027f: data_buf = 8'h53;
			13'h0280: data_buf = 8'h43;
			13'h0281: data_buf = 8'hc3;
			13'h0282: data_buf = 8'h48;
			13'h0283: data_buf = 8'h52;
			13'h0284: data_buf = 8'h24;
			13'h0285: data_buf = 8'hc8;
			13'h0286: data_buf = 8'h45;
			13'h0287: data_buf = 8'h58;
			13'h0288: data_buf = 8'h24;
			13'h0289: data_buf = 8'hc2;
			13'h028a: data_buf = 8'h49;
			13'h028b: data_buf = 8'h4e;
			13'h028c: data_buf = 8'h24;
			13'h028d: data_buf = 8'hcc;
			13'h028e: data_buf = 8'h45;
			13'h028f: data_buf = 8'h46;
			13'h0290: data_buf = 8'h54;
			13'h0291: data_buf = 8'h24;
			13'h0292: data_buf = 8'hd2;
			13'h0293: data_buf = 8'h49;
			13'h0294: data_buf = 8'h47;
			13'h0295: data_buf = 8'h48;
			13'h0296: data_buf = 8'h54;
			13'h0297: data_buf = 8'h24;
			13'h0298: data_buf = 8'hcd;
			13'h0299: data_buf = 8'h49;
			13'h029a: data_buf = 8'h44;
			13'h029b: data_buf = 8'h24;
			13'h029c: data_buf = 8'h80;
			13'h029d: data_buf = 8'h97;
			13'h029e: data_buf = 8'h08;
			13'h029f: data_buf = 8'h94;
			13'h02a0: data_buf = 8'h07;
			13'h02a1: data_buf = 8'h6f;
			13'h02a2: data_buf = 8'h0c;
			13'h02a3: data_buf = 8'he4;
			13'h02a4: data_buf = 8'h09;
			13'h02a5: data_buf = 8'h76;
			13'h02a6: data_buf = 8'h0b;
			13'h02a7: data_buf = 8'hab;
			13'h02a8: data_buf = 8'h0e;
			13'h02a9: data_buf = 8'ha5;
			13'h02aa: data_buf = 8'h0b;
			13'h02ab: data_buf = 8'hfb;
			13'h02ac: data_buf = 8'h09;
			13'h02ad: data_buf = 8'ha1;
			13'h02ae: data_buf = 8'h09;
			13'h02af: data_buf = 8'h84;
			13'h02b0: data_buf = 8'h09;
			13'h02b1: data_buf = 8'h73;
			13'h02b2: data_buf = 8'h0a;
			13'h02b3: data_buf = 8'h5d;
			13'h02b4: data_buf = 8'h08;
			13'h02b5: data_buf = 8'h90;
			13'h02b6: data_buf = 8'h09;
			13'h02b7: data_buf = 8'hbf;
			13'h02b8: data_buf = 8'h09;
			13'h02b9: data_buf = 8'he6;
			13'h02ba: data_buf = 8'h09;
			13'h02bb: data_buf = 8'h95;
			13'h02bc: data_buf = 8'h08;
			13'h02bd: data_buf = 8'he4;
			13'h02be: data_buf = 8'h13;
			13'h02bf: data_buf = 8'h55;
			13'h02c0: data_buf = 8'h0a;
			13'h02c1: data_buf = 8'hd6;
			13'h02c2: data_buf = 8'h08;
			13'h02c3: data_buf = 8'hea;
			13'h02c4: data_buf = 8'h13;
			13'h02c5: data_buf = 8'h89;
			13'h02c6: data_buf = 8'h10;
			13'h02c7: data_buf = 8'h33;
			13'h02c8: data_buf = 8'h14;
			13'h02c9: data_buf = 8'h7b;
			13'h02ca: data_buf = 8'h1b;
			13'h02cb: data_buf = 8'he6;
			13'h02cc: data_buf = 8'h09;
			13'h02cd: data_buf = 8'h61;
			13'h02ce: data_buf = 8'h1b;
			13'h02cf: data_buf = 8'h54;
			13'h02d0: data_buf = 8'h1b;
			13'h02d1: data_buf = 8'h59;
			13'h02d2: data_buf = 8'h1b;
			13'h02d3: data_buf = 8'h8d;
			13'h02d4: data_buf = 8'h1c;
			13'h02d5: data_buf = 8'h99;
			13'h02d6: data_buf = 8'h80;
			13'h02d7: data_buf = 8'h9c;
			13'h02d8: data_buf = 8'h80;
			13'h02d9: data_buf = 8'h97;
			13'h02da: data_buf = 8'h0a;
			13'h02db: data_buf = 8'hc3;
			13'h02dc: data_buf = 8'h08;
			13'h02dd: data_buf = 8'h09;
			13'h02de: data_buf = 8'h07;
			13'h02df: data_buf = 8'h3e;
			13'h02e0: data_buf = 8'h09;
			13'h02e1: data_buf = 8'he6;
			13'h02e2: data_buf = 8'h09;
			13'h02e3: data_buf = 8'he6;
			13'h02e4: data_buf = 8'h09;
			13'h02e5: data_buf = 8'h01;
			13'h02e6: data_buf = 8'h05;
			13'h02e7: data_buf = 8'h79;
			13'h02e8: data_buf = 8'h1d;
			13'h02e9: data_buf = 8'h18;
			13'h02ea: data_buf = 8'h79;
			13'h02eb: data_buf = 8'h51;
			13'h02ec: data_buf = 8'h14;
			13'h02ed: data_buf = 8'h7c;
			13'h02ee: data_buf = 8'h8f;
			13'h02ef: data_buf = 8'h15;
			13'h02f0: data_buf = 8'h7c;
			13'h02f1: data_buf = 8'hf0;
			13'h02f2: data_buf = 8'h15;
			13'h02f3: data_buf = 8'h7f;
			13'h02f4: data_buf = 8'h3e;
			13'h02f5: data_buf = 8'h19;
			13'h02f6: data_buf = 8'h50;
			13'h02f7: data_buf = 8'h04;
			13'h02f8: data_buf = 8'h0e;
			13'h02f9: data_buf = 8'h46;
			13'h02fa: data_buf = 8'h03;
			13'h02fb: data_buf = 8'h0e;
			13'h02fc: data_buf = 8'h4e;
			13'h02fd: data_buf = 8'h46;
			13'h02fe: data_buf = 8'h53;
			13'h02ff: data_buf = 8'h4e;
			13'h0300: data_buf = 8'h52;
			13'h0301: data_buf = 8'h47;
			13'h0302: data_buf = 8'h4f;
			13'h0303: data_buf = 8'h44;
			13'h0304: data_buf = 8'h46;
			13'h0305: data_buf = 8'h43;
			13'h0306: data_buf = 8'h4f;
			13'h0307: data_buf = 8'h56;
			13'h0308: data_buf = 8'h4f;
			13'h0309: data_buf = 8'h4d;
			13'h030a: data_buf = 8'h55;
			13'h030b: data_buf = 8'h4c;
			13'h030c: data_buf = 8'h42;
			13'h030d: data_buf = 8'h53;
			13'h030e: data_buf = 8'h44;
			13'h030f: data_buf = 8'h44;
			13'h0310: data_buf = 8'h2f;
			13'h0311: data_buf = 8'h30;
			13'h0312: data_buf = 8'h49;
			13'h0313: data_buf = 8'h44;
			13'h0314: data_buf = 8'h54;
			13'h0315: data_buf = 8'h4d;
			13'h0316: data_buf = 8'h4f;
			13'h0317: data_buf = 8'h53;
			13'h0318: data_buf = 8'h4c;
			13'h0319: data_buf = 8'h53;
			13'h031a: data_buf = 8'h53;
			13'h031b: data_buf = 8'h54;
			13'h031c: data_buf = 8'h43;
			13'h031d: data_buf = 8'h4e;
			13'h031e: data_buf = 8'h55;
			13'h031f: data_buf = 8'h46;
			13'h0320: data_buf = 8'h4d;
			13'h0321: data_buf = 8'h4f;
			13'h0322: data_buf = 8'h48;
			13'h0323: data_buf = 8'h58;
			13'h0324: data_buf = 8'h42;
			13'h0325: data_buf = 8'h4e;
			13'h0326: data_buf = 8'hc3;
			13'h0327: data_buf = 8'hbc;
			13'h0328: data_buf = 8'h00;
			13'h0329: data_buf = 8'hc3;
			13'h032a: data_buf = 8'h14;
			13'h032b: data_buf = 8'h09;
			13'h032c: data_buf = 8'hd3;
			13'h032d: data_buf = 8'h00;
			13'h032e: data_buf = 8'hc9;
			13'h032f: data_buf = 8'hd6;
			13'h0330: data_buf = 8'h00;
			13'h0331: data_buf = 8'h6f;
			13'h0332: data_buf = 8'h7c;
			13'h0333: data_buf = 8'hde;
			13'h0334: data_buf = 8'h00;
			13'h0335: data_buf = 8'h67;
			13'h0336: data_buf = 8'h78;
			13'h0337: data_buf = 8'hde;
			13'h0338: data_buf = 8'h00;
			13'h0339: data_buf = 8'h47;
			13'h033a: data_buf = 8'h3e;
			13'h033b: data_buf = 8'h00;
			13'h033c: data_buf = 8'hc9;
			13'h033d: data_buf = 8'h00;
			13'h033e: data_buf = 8'h00;
			13'h033f: data_buf = 8'h00;
			13'h0340: data_buf = 8'h35;
			13'h0341: data_buf = 8'h4a;
			13'h0342: data_buf = 8'hca;
			13'h0343: data_buf = 8'h99;
			13'h0344: data_buf = 8'h39;
			13'h0345: data_buf = 8'h1c;
			13'h0346: data_buf = 8'h76;
			13'h0347: data_buf = 8'h98;
			13'h0348: data_buf = 8'h22;
			13'h0349: data_buf = 8'h95;
			13'h034a: data_buf = 8'hb3;
			13'h034b: data_buf = 8'h98;
			13'h034c: data_buf = 8'h0a;
			13'h034d: data_buf = 8'hdd;
			13'h034e: data_buf = 8'h47;
			13'h034f: data_buf = 8'h98;
			13'h0350: data_buf = 8'h53;
			13'h0351: data_buf = 8'hd1;
			13'h0352: data_buf = 8'h99;
			13'h0353: data_buf = 8'h99;
			13'h0354: data_buf = 8'h0a;
			13'h0355: data_buf = 8'h1a;
			13'h0356: data_buf = 8'h9f;
			13'h0357: data_buf = 8'h98;
			13'h0358: data_buf = 8'h65;
			13'h0359: data_buf = 8'hbc;
			13'h035a: data_buf = 8'hcd;
			13'h035b: data_buf = 8'h98;
			13'h035c: data_buf = 8'hd6;
			13'h035d: data_buf = 8'h77;
			13'h035e: data_buf = 8'h3e;
			13'h035f: data_buf = 8'h98;
			13'h0360: data_buf = 8'h52;
			13'h0361: data_buf = 8'hc7;
			13'h0362: data_buf = 8'h4f;
			13'h0363: data_buf = 8'h80;
			13'h0364: data_buf = 8'hdb;
			13'h0365: data_buf = 8'h00;
			13'h0366: data_buf = 8'hc9;
			13'h0367: data_buf = 8'h01;
			13'h0368: data_buf = 8'hff;
			13'h0369: data_buf = 8'h1c;
			13'h036a: data_buf = 8'h00;
			13'h036b: data_buf = 8'h00;
			13'h036c: data_buf = 8'h14;
			13'h036d: data_buf = 8'h00;
			13'h036e: data_buf = 8'h14;
			13'h036f: data_buf = 8'h00;
			13'h0370: data_buf = 8'h00;
			13'h0371: data_buf = 8'h00;
			13'h0372: data_buf = 8'h00;
			13'h0373: data_buf = 8'h00;
			13'h0374: data_buf = 8'hc3;
			13'h0375: data_buf = 8'h3a;
			13'h0376: data_buf = 8'h06;
			13'h0377: data_buf = 8'hc3;
			13'h0378: data_buf = 8'h00;
			13'h0379: data_buf = 8'h00;
			13'h037a: data_buf = 8'hc3;
			13'h037b: data_buf = 8'h00;
			13'h037c: data_buf = 8'h00;
			13'h037d: data_buf = 8'hc3;
			13'h037e: data_buf = 8'h00;
			13'h037f: data_buf = 8'h00;
			13'h0380: data_buf = 8'ha2;
			13'h0381: data_buf = 8'h81;
			13'h0382: data_buf = 8'hfe;
			13'h0383: data_buf = 8'hff;
			13'h0384: data_buf = 8'h3f;
			13'h0385: data_buf = 8'h81;
			13'h0386: data_buf = 8'h20;
			13'h0387: data_buf = 8'h45;
			13'h0388: data_buf = 8'h72;
			13'h0389: data_buf = 8'h72;
			13'h038a: data_buf = 8'h6f;
			13'h038b: data_buf = 8'h72;
			13'h038c: data_buf = 8'h00;
			13'h038d: data_buf = 8'h20;
			13'h038e: data_buf = 8'h69;
			13'h038f: data_buf = 8'h6e;
			13'h0390: data_buf = 8'h20;
			13'h0391: data_buf = 8'h00;
			13'h0392: data_buf = 8'h4f;
			13'h0393: data_buf = 8'h6b;
			13'h0394: data_buf = 8'h0d;
			13'h0395: data_buf = 8'h0a;
			13'h0396: data_buf = 8'h00;
			13'h0397: data_buf = 8'h00;
			13'h0398: data_buf = 8'h42;
			13'h0399: data_buf = 8'h72;
			13'h039a: data_buf = 8'h65;
			13'h039b: data_buf = 8'h61;
			13'h039c: data_buf = 8'h6b;
			13'h039d: data_buf = 8'h00;
			13'h039e: data_buf = 8'h21;
			13'h039f: data_buf = 8'h04;
			13'h03a0: data_buf = 8'h00;
			13'h03a1: data_buf = 8'h39;
			13'h03a2: data_buf = 8'h7e;
			13'h03a3: data_buf = 8'h23;
			13'h03a4: data_buf = 8'hfe;
			13'h03a5: data_buf = 8'h81;
			13'h03a6: data_buf = 8'hc0;
			13'h03a7: data_buf = 8'h4e;
			13'h03a8: data_buf = 8'h23;
			13'h03a9: data_buf = 8'h46;
			13'h03aa: data_buf = 8'h23;
			13'h03ab: data_buf = 8'he5;
			13'h03ac: data_buf = 8'h69;
			13'h03ad: data_buf = 8'h60;
			13'h03ae: data_buf = 8'h7a;
			13'h03af: data_buf = 8'hb3;
			13'h03b0: data_buf = 8'heb;
			13'h03b1: data_buf = 8'hca;
			13'h03b2: data_buf = 8'hb8;
			13'h03b3: data_buf = 8'h03;
			13'h03b4: data_buf = 8'heb;
			13'h03b5: data_buf = 8'hcd;
			13'h03b6: data_buf = 8'hbd;
			13'h03b7: data_buf = 8'h06;
			13'h03b8: data_buf = 8'h01;
			13'h03b9: data_buf = 8'h0d;
			13'h03ba: data_buf = 8'h00;
			13'h03bb: data_buf = 8'he1;
			13'h03bc: data_buf = 8'hc8;
			13'h03bd: data_buf = 8'h09;
			13'h03be: data_buf = 8'hc3;
			13'h03bf: data_buf = 8'ha2;
			13'h03c0: data_buf = 8'h03;
			13'h03c1: data_buf = 8'hcd;
			13'h03c2: data_buf = 8'hdb;
			13'h03c3: data_buf = 8'h03;
			13'h03c4: data_buf = 8'hc5;
			13'h03c5: data_buf = 8'he3;
			13'h03c6: data_buf = 8'hc1;
			13'h03c7: data_buf = 8'hcd;
			13'h03c8: data_buf = 8'hbd;
			13'h03c9: data_buf = 8'h06;
			13'h03ca: data_buf = 8'h7e;
			13'h03cb: data_buf = 8'h02;
			13'h03cc: data_buf = 8'hc8;
			13'h03cd: data_buf = 8'h0b;
			13'h03ce: data_buf = 8'h2b;
			13'h03cf: data_buf = 8'hc3;
			13'h03d0: data_buf = 8'hc7;
			13'h03d1: data_buf = 8'h03;
			13'h03d2: data_buf = 8'he5;
			13'h03d3: data_buf = 8'h2a;
			13'h03d4: data_buf = 8'h1f;
			13'h03d5: data_buf = 8'h81;
			13'h03d6: data_buf = 8'h06;
			13'h03d7: data_buf = 8'h00;
			13'h03d8: data_buf = 8'h09;
			13'h03d9: data_buf = 8'h09;
			13'h03da: data_buf = 8'h3e;
			13'h03db: data_buf = 8'he5;
			13'h03dc: data_buf = 8'h3e;
			13'h03dd: data_buf = 8'hd0;
			13'h03de: data_buf = 8'h95;
			13'h03df: data_buf = 8'h6f;
			13'h03e0: data_buf = 8'h3e;
			13'h03e1: data_buf = 8'hff;
			13'h03e2: data_buf = 8'h9c;
			13'h03e3: data_buf = 8'hda;
			13'h03e4: data_buf = 8'hea;
			13'h03e5: data_buf = 8'h03;
			13'h03e6: data_buf = 8'h67;
			13'h03e7: data_buf = 8'h39;
			13'h03e8: data_buf = 8'he1;
			13'h03e9: data_buf = 8'hd8;
			13'h03ea: data_buf = 8'h1e;
			13'h03eb: data_buf = 8'h0c;
			13'h03ec: data_buf = 8'hc3;
			13'h03ed: data_buf = 8'h09;
			13'h03ee: data_buf = 8'h04;
			13'h03ef: data_buf = 8'h2a;
			13'h03f0: data_buf = 8'h0e;
			13'h03f1: data_buf = 8'h81;
			13'h03f2: data_buf = 8'h22;
			13'h03f3: data_buf = 8'ha1;
			13'h03f4: data_buf = 8'h80;
			13'h03f5: data_buf = 8'h1e;
			13'h03f6: data_buf = 8'h02;
			13'h03f7: data_buf = 8'h01;
			13'h03f8: data_buf = 8'h1e;
			13'h03f9: data_buf = 8'h14;
			13'h03fa: data_buf = 8'h01;
			13'h03fb: data_buf = 8'h1e;
			13'h03fc: data_buf = 8'h00;
			13'h03fd: data_buf = 8'h01;
			13'h03fe: data_buf = 8'h1e;
			13'h03ff: data_buf = 8'h12;
			13'h0400: data_buf = 8'h01;
			13'h0401: data_buf = 8'h1e;
			13'h0402: data_buf = 8'h22;
			13'h0403: data_buf = 8'h01;
			13'h0404: data_buf = 8'h1e;
			13'h0405: data_buf = 8'h0a;
			13'h0406: data_buf = 8'h01;
			13'h0407: data_buf = 8'h1e;
			13'h0408: data_buf = 8'h18;
			13'h0409: data_buf = 8'hcd;
			13'h040a: data_buf = 8'h27;
			13'h040b: data_buf = 8'h05;
			13'h040c: data_buf = 8'h32;
			13'h040d: data_buf = 8'h8a;
			13'h040e: data_buf = 8'h80;
			13'h040f: data_buf = 8'hcd;
			13'h0410: data_buf = 8'he8;
			13'h0411: data_buf = 8'h0a;
			13'h0412: data_buf = 8'h21;
			13'h0413: data_buf = 8'hfc;
			13'h0414: data_buf = 8'h02;
			13'h0415: data_buf = 8'h57;
			13'h0416: data_buf = 8'h3e;
			13'h0417: data_buf = 8'h3f;
			13'h0418: data_buf = 8'hcd;
			13'h0419: data_buf = 8'hce;
			13'h041a: data_buf = 8'h06;
			13'h041b: data_buf = 8'h19;
			13'h041c: data_buf = 8'h7e;
			13'h041d: data_buf = 8'hcd;
			13'h041e: data_buf = 8'hce;
			13'h041f: data_buf = 8'h06;
			13'h0420: data_buf = 8'hcd;
			13'h0421: data_buf = 8'h4d;
			13'h0422: data_buf = 8'h08;
			13'h0423: data_buf = 8'hcd;
			13'h0424: data_buf = 8'hce;
			13'h0425: data_buf = 8'h06;
			13'h0426: data_buf = 8'h21;
			13'h0427: data_buf = 8'h86;
			13'h0428: data_buf = 8'h03;
			13'h0429: data_buf = 8'hcd;
			13'h042a: data_buf = 8'h93;
			13'h042b: data_buf = 8'h11;
			13'h042c: data_buf = 8'h2a;
			13'h042d: data_buf = 8'ha1;
			13'h042e: data_buf = 8'h80;
			13'h042f: data_buf = 8'h11;
			13'h0430: data_buf = 8'hfe;
			13'h0431: data_buf = 8'hff;
			13'h0432: data_buf = 8'hcd;
			13'h0433: data_buf = 8'hbd;
			13'h0434: data_buf = 8'h06;
			13'h0435: data_buf = 8'hca;
			13'h0436: data_buf = 8'h4e;
			13'h0437: data_buf = 8'h00;
			13'h0438: data_buf = 8'h7c;
			13'h0439: data_buf = 8'ha5;
			13'h043a: data_buf = 8'h3c;
			13'h043b: data_buf = 8'hc4;
			13'h043c: data_buf = 8'h2e;
			13'h043d: data_buf = 8'h18;
			13'h043e: data_buf = 8'h3e;
			13'h043f: data_buf = 8'hc1;
			13'h0440: data_buf = 8'haf;
			13'h0441: data_buf = 8'h32;
			13'h0442: data_buf = 8'h8a;
			13'h0443: data_buf = 8'h80;
			13'h0444: data_buf = 8'hcd;
			13'h0445: data_buf = 8'he8;
			13'h0446: data_buf = 8'h0a;
			13'h0447: data_buf = 8'h21;
			13'h0448: data_buf = 8'h92;
			13'h0449: data_buf = 8'h03;
			13'h044a: data_buf = 8'hcd;
			13'h044b: data_buf = 8'h93;
			13'h044c: data_buf = 8'h11;
			13'h044d: data_buf = 8'h21;
			13'h044e: data_buf = 8'hff;
			13'h044f: data_buf = 8'hff;
			13'h0450: data_buf = 8'h22;
			13'h0451: data_buf = 8'ha1;
			13'h0452: data_buf = 8'h80;
			13'h0453: data_buf = 8'hcd;
			13'h0454: data_buf = 8'h3a;
			13'h0455: data_buf = 8'h06;
			13'h0456: data_buf = 8'hda;
			13'h0457: data_buf = 8'h4d;
			13'h0458: data_buf = 8'h04;
			13'h0459: data_buf = 8'hcd;
			13'h045a: data_buf = 8'h4d;
			13'h045b: data_buf = 8'h08;
			13'h045c: data_buf = 8'h3c;
			13'h045d: data_buf = 8'h3d;
			13'h045e: data_buf = 8'hca;
			13'h045f: data_buf = 8'h4d;
			13'h0460: data_buf = 8'h04;
			13'h0461: data_buf = 8'hf5;
			13'h0462: data_buf = 8'hcd;
			13'h0463: data_buf = 8'h19;
			13'h0464: data_buf = 8'h09;
			13'h0465: data_buf = 8'hd5;
			13'h0466: data_buf = 8'hcd;
			13'h0467: data_buf = 8'h51;
			13'h0468: data_buf = 8'h05;
			13'h0469: data_buf = 8'h47;
			13'h046a: data_buf = 8'hd1;
			13'h046b: data_buf = 8'hf1;
			13'h046c: data_buf = 8'hd2;
			13'h046d: data_buf = 8'h2d;
			13'h046e: data_buf = 8'h08;
			13'h046f: data_buf = 8'hd5;
			13'h0470: data_buf = 8'hc5;
			13'h0471: data_buf = 8'haf;
			13'h0472: data_buf = 8'h32;
			13'h0473: data_buf = 8'h11;
			13'h0474: data_buf = 8'h81;
			13'h0475: data_buf = 8'hcd;
			13'h0476: data_buf = 8'h4d;
			13'h0477: data_buf = 8'h08;
			13'h0478: data_buf = 8'hb7;
			13'h0479: data_buf = 8'hf5;
			13'h047a: data_buf = 8'hcd;
			13'h047b: data_buf = 8'he1;
			13'h047c: data_buf = 8'h04;
			13'h047d: data_buf = 8'hda;
			13'h047e: data_buf = 8'h86;
			13'h047f: data_buf = 8'h04;
			13'h0480: data_buf = 8'hf1;
			13'h0481: data_buf = 8'hf5;
			13'h0482: data_buf = 8'hca;
			13'h0483: data_buf = 8'hba;
			13'h0484: data_buf = 8'h09;
			13'h0485: data_buf = 8'hb7;
			13'h0486: data_buf = 8'hc5;
			13'h0487: data_buf = 8'hd2;
			13'h0488: data_buf = 8'h9d;
			13'h0489: data_buf = 8'h04;
			13'h048a: data_buf = 8'heb;
			13'h048b: data_buf = 8'h2a;
			13'h048c: data_buf = 8'h1b;
			13'h048d: data_buf = 8'h81;
			13'h048e: data_buf = 8'h1a;
			13'h048f: data_buf = 8'h02;
			13'h0490: data_buf = 8'h03;
			13'h0491: data_buf = 8'h13;
			13'h0492: data_buf = 8'hcd;
			13'h0493: data_buf = 8'hbd;
			13'h0494: data_buf = 8'h06;
			13'h0495: data_buf = 8'hc2;
			13'h0496: data_buf = 8'h8e;
			13'h0497: data_buf = 8'h04;
			13'h0498: data_buf = 8'h60;
			13'h0499: data_buf = 8'h69;
			13'h049a: data_buf = 8'h22;
			13'h049b: data_buf = 8'h1b;
			13'h049c: data_buf = 8'h81;
			13'h049d: data_buf = 8'hd1;
			13'h049e: data_buf = 8'hf1;
			13'h049f: data_buf = 8'hca;
			13'h04a0: data_buf = 8'hc4;
			13'h04a1: data_buf = 8'h04;
			13'h04a2: data_buf = 8'h2a;
			13'h04a3: data_buf = 8'h1b;
			13'h04a4: data_buf = 8'h81;
			13'h04a5: data_buf = 8'he3;
			13'h04a6: data_buf = 8'hc1;
			13'h04a7: data_buf = 8'h09;
			13'h04a8: data_buf = 8'he5;
			13'h04a9: data_buf = 8'hcd;
			13'h04aa: data_buf = 8'hc1;
			13'h04ab: data_buf = 8'h03;
			13'h04ac: data_buf = 8'he1;
			13'h04ad: data_buf = 8'h22;
			13'h04ae: data_buf = 8'h1b;
			13'h04af: data_buf = 8'h81;
			13'h04b0: data_buf = 8'heb;
			13'h04b1: data_buf = 8'h74;
			13'h04b2: data_buf = 8'hd1;
			13'h04b3: data_buf = 8'h23;
			13'h04b4: data_buf = 8'h23;
			13'h04b5: data_buf = 8'h73;
			13'h04b6: data_buf = 8'h23;
			13'h04b7: data_buf = 8'h72;
			13'h04b8: data_buf = 8'h23;
			13'h04b9: data_buf = 8'h11;
			13'h04ba: data_buf = 8'ha6;
			13'h04bb: data_buf = 8'h80;
			13'h04bc: data_buf = 8'h1a;
			13'h04bd: data_buf = 8'h77;
			13'h04be: data_buf = 8'h23;
			13'h04bf: data_buf = 8'h13;
			13'h04c0: data_buf = 8'hb7;
			13'h04c1: data_buf = 8'hc2;
			13'h04c2: data_buf = 8'hbc;
			13'h04c3: data_buf = 8'h04;
			13'h04c4: data_buf = 8'hcd;
			13'h04c5: data_buf = 8'h0d;
			13'h04c6: data_buf = 8'h05;
			13'h04c7: data_buf = 8'h23;
			13'h04c8: data_buf = 8'heb;
			13'h04c9: data_buf = 8'h62;
			13'h04ca: data_buf = 8'h6b;
			13'h04cb: data_buf = 8'h7e;
			13'h04cc: data_buf = 8'h23;
			13'h04cd: data_buf = 8'hb6;
			13'h04ce: data_buf = 8'hca;
			13'h04cf: data_buf = 8'h4d;
			13'h04d0: data_buf = 8'h04;
			13'h04d1: data_buf = 8'h23;
			13'h04d2: data_buf = 8'h23;
			13'h04d3: data_buf = 8'h23;
			13'h04d4: data_buf = 8'haf;
			13'h04d5: data_buf = 8'hbe;
			13'h04d6: data_buf = 8'h23;
			13'h04d7: data_buf = 8'hc2;
			13'h04d8: data_buf = 8'hd5;
			13'h04d9: data_buf = 8'h04;
			13'h04da: data_buf = 8'heb;
			13'h04db: data_buf = 8'h73;
			13'h04dc: data_buf = 8'h23;
			13'h04dd: data_buf = 8'h72;
			13'h04de: data_buf = 8'hc3;
			13'h04df: data_buf = 8'hc9;
			13'h04e0: data_buf = 8'h04;
			13'h04e1: data_buf = 8'h2a;
			13'h04e2: data_buf = 8'ha3;
			13'h04e3: data_buf = 8'h80;
			13'h04e4: data_buf = 8'h44;
			13'h04e5: data_buf = 8'h4d;
			13'h04e6: data_buf = 8'h7e;
			13'h04e7: data_buf = 8'h23;
			13'h04e8: data_buf = 8'hb6;
			13'h04e9: data_buf = 8'h2b;
			13'h04ea: data_buf = 8'hc8;
			13'h04eb: data_buf = 8'h23;
			13'h04ec: data_buf = 8'h23;
			13'h04ed: data_buf = 8'h7e;
			13'h04ee: data_buf = 8'h23;
			13'h04ef: data_buf = 8'h66;
			13'h04f0: data_buf = 8'h6f;
			13'h04f1: data_buf = 8'hcd;
			13'h04f2: data_buf = 8'hbd;
			13'h04f3: data_buf = 8'h06;
			13'h04f4: data_buf = 8'h60;
			13'h04f5: data_buf = 8'h69;
			13'h04f6: data_buf = 8'h7e;
			13'h04f7: data_buf = 8'h23;
			13'h04f8: data_buf = 8'h66;
			13'h04f9: data_buf = 8'h6f;
			13'h04fa: data_buf = 8'h3f;
			13'h04fb: data_buf = 8'hc8;
			13'h04fc: data_buf = 8'h3f;
			13'h04fd: data_buf = 8'hd0;
			13'h04fe: data_buf = 8'hc3;
			13'h04ff: data_buf = 8'he4;
			13'h0500: data_buf = 8'h04;
			13'h0501: data_buf = 8'hc0;
			13'h0502: data_buf = 8'h2a;
			13'h0503: data_buf = 8'ha3;
			13'h0504: data_buf = 8'h80;
			13'h0505: data_buf = 8'haf;
			13'h0506: data_buf = 8'h77;
			13'h0507: data_buf = 8'h23;
			13'h0508: data_buf = 8'h77;
			13'h0509: data_buf = 8'h23;
			13'h050a: data_buf = 8'h22;
			13'h050b: data_buf = 8'h1b;
			13'h050c: data_buf = 8'h81;
			13'h050d: data_buf = 8'h2a;
			13'h050e: data_buf = 8'ha3;
			13'h050f: data_buf = 8'h80;
			13'h0510: data_buf = 8'h2b;
			13'h0511: data_buf = 8'h22;
			13'h0512: data_buf = 8'h13;
			13'h0513: data_buf = 8'h81;
			13'h0514: data_buf = 8'h2a;
			13'h0515: data_buf = 8'hf4;
			13'h0516: data_buf = 8'h80;
			13'h0517: data_buf = 8'h22;
			13'h0518: data_buf = 8'h08;
			13'h0519: data_buf = 8'h81;
			13'h051a: data_buf = 8'haf;
			13'h051b: data_buf = 8'hcd;
			13'h051c: data_buf = 8'h5d;
			13'h051d: data_buf = 8'h08;
			13'h051e: data_buf = 8'h2a;
			13'h051f: data_buf = 8'h1b;
			13'h0520: data_buf = 8'h81;
			13'h0521: data_buf = 8'h22;
			13'h0522: data_buf = 8'h1d;
			13'h0523: data_buf = 8'h81;
			13'h0524: data_buf = 8'h22;
			13'h0525: data_buf = 8'h1f;
			13'h0526: data_buf = 8'h81;
			13'h0527: data_buf = 8'hc1;
			13'h0528: data_buf = 8'h2a;
			13'h0529: data_buf = 8'h9f;
			13'h052a: data_buf = 8'h80;
			13'h052b: data_buf = 8'hf9;
			13'h052c: data_buf = 8'h21;
			13'h052d: data_buf = 8'hf8;
			13'h052e: data_buf = 8'h80;
			13'h052f: data_buf = 8'h22;
			13'h0530: data_buf = 8'hf6;
			13'h0531: data_buf = 8'h80;
			13'h0532: data_buf = 8'haf;
			13'h0533: data_buf = 8'h6f;
			13'h0534: data_buf = 8'h67;
			13'h0535: data_buf = 8'h22;
			13'h0536: data_buf = 8'h19;
			13'h0537: data_buf = 8'h81;
			13'h0538: data_buf = 8'h32;
			13'h0539: data_buf = 8'h10;
			13'h053a: data_buf = 8'h81;
			13'h053b: data_buf = 8'h22;
			13'h053c: data_buf = 8'h23;
			13'h053d: data_buf = 8'h81;
			13'h053e: data_buf = 8'he5;
			13'h053f: data_buf = 8'hc5;
			13'h0540: data_buf = 8'h2a;
			13'h0541: data_buf = 8'h13;
			13'h0542: data_buf = 8'h81;
			13'h0543: data_buf = 8'hc9;
			13'h0544: data_buf = 8'h3e;
			13'h0545: data_buf = 8'h3f;
			13'h0546: data_buf = 8'hcd;
			13'h0547: data_buf = 8'hce;
			13'h0548: data_buf = 8'h06;
			13'h0549: data_buf = 8'h3e;
			13'h054a: data_buf = 8'h20;
			13'h054b: data_buf = 8'hcd;
			13'h054c: data_buf = 8'hce;
			13'h054d: data_buf = 8'h06;
			13'h054e: data_buf = 8'hc3;
			13'h054f: data_buf = 8'h93;
			13'h0550: data_buf = 8'h80;
			13'h0551: data_buf = 8'haf;
			13'h0552: data_buf = 8'h32;
			13'h0553: data_buf = 8'hf3;
			13'h0554: data_buf = 8'h80;
			13'h0555: data_buf = 8'h0e;
			13'h0556: data_buf = 8'h05;
			13'h0557: data_buf = 8'h11;
			13'h0558: data_buf = 8'ha6;
			13'h0559: data_buf = 8'h80;
			13'h055a: data_buf = 8'h7e;
			13'h055b: data_buf = 8'hfe;
			13'h055c: data_buf = 8'h20;
			13'h055d: data_buf = 8'hca;
			13'h055e: data_buf = 8'hd9;
			13'h055f: data_buf = 8'h05;
			13'h0560: data_buf = 8'h47;
			13'h0561: data_buf = 8'hfe;
			13'h0562: data_buf = 8'h22;
			13'h0563: data_buf = 8'hca;
			13'h0564: data_buf = 8'hf9;
			13'h0565: data_buf = 8'h05;
			13'h0566: data_buf = 8'hb7;
			13'h0567: data_buf = 8'hca;
			13'h0568: data_buf = 8'h00;
			13'h0569: data_buf = 8'h06;
			13'h056a: data_buf = 8'h3a;
			13'h056b: data_buf = 8'hf3;
			13'h056c: data_buf = 8'h80;
			13'h056d: data_buf = 8'hb7;
			13'h056e: data_buf = 8'h7e;
			13'h056f: data_buf = 8'hc2;
			13'h0570: data_buf = 8'hd9;
			13'h0571: data_buf = 8'h05;
			13'h0572: data_buf = 8'hfe;
			13'h0573: data_buf = 8'h3f;
			13'h0574: data_buf = 8'h3e;
			13'h0575: data_buf = 8'h9e;
			13'h0576: data_buf = 8'hca;
			13'h0577: data_buf = 8'hd9;
			13'h0578: data_buf = 8'h05;
			13'h0579: data_buf = 8'h7e;
			13'h057a: data_buf = 8'hfe;
			13'h057b: data_buf = 8'h30;
			13'h057c: data_buf = 8'hda;
			13'h057d: data_buf = 8'h84;
			13'h057e: data_buf = 8'h05;
			13'h057f: data_buf = 8'hfe;
			13'h0580: data_buf = 8'h3c;
			13'h0581: data_buf = 8'hda;
			13'h0582: data_buf = 8'hd9;
			13'h0583: data_buf = 8'h05;
			13'h0584: data_buf = 8'hd5;
			13'h0585: data_buf = 8'h11;
			13'h0586: data_buf = 8'h7d;
			13'h0587: data_buf = 8'h01;
			13'h0588: data_buf = 8'hc5;
			13'h0589: data_buf = 8'h01;
			13'h058a: data_buf = 8'hd5;
			13'h058b: data_buf = 8'h05;
			13'h058c: data_buf = 8'hc5;
			13'h058d: data_buf = 8'h06;
			13'h058e: data_buf = 8'h7f;
			13'h058f: data_buf = 8'h7e;
			13'h0590: data_buf = 8'hfe;
			13'h0591: data_buf = 8'h61;
			13'h0592: data_buf = 8'hda;
			13'h0593: data_buf = 8'h9d;
			13'h0594: data_buf = 8'h05;
			13'h0595: data_buf = 8'hfe;
			13'h0596: data_buf = 8'h7b;
			13'h0597: data_buf = 8'hd2;
			13'h0598: data_buf = 8'h9d;
			13'h0599: data_buf = 8'h05;
			13'h059a: data_buf = 8'he6;
			13'h059b: data_buf = 8'h5f;
			13'h059c: data_buf = 8'h77;
			13'h059d: data_buf = 8'h4e;
			13'h059e: data_buf = 8'heb;
			13'h059f: data_buf = 8'h23;
			13'h05a0: data_buf = 8'hb6;
			13'h05a1: data_buf = 8'hf2;
			13'h05a2: data_buf = 8'h9f;
			13'h05a3: data_buf = 8'h05;
			13'h05a4: data_buf = 8'h04;
			13'h05a5: data_buf = 8'h7e;
			13'h05a6: data_buf = 8'he6;
			13'h05a7: data_buf = 8'h7f;
			13'h05a8: data_buf = 8'hc8;
			13'h05a9: data_buf = 8'hb9;
			13'h05aa: data_buf = 8'hc2;
			13'h05ab: data_buf = 8'h9f;
			13'h05ac: data_buf = 8'h05;
			13'h05ad: data_buf = 8'heb;
			13'h05ae: data_buf = 8'he5;
			13'h05af: data_buf = 8'h13;
			13'h05b0: data_buf = 8'h1a;
			13'h05b1: data_buf = 8'hb7;
			13'h05b2: data_buf = 8'hfa;
			13'h05b3: data_buf = 8'hd1;
			13'h05b4: data_buf = 8'h05;
			13'h05b5: data_buf = 8'h4f;
			13'h05b6: data_buf = 8'h78;
			13'h05b7: data_buf = 8'hfe;
			13'h05b8: data_buf = 8'h88;
			13'h05b9: data_buf = 8'hc2;
			13'h05ba: data_buf = 8'hc0;
			13'h05bb: data_buf = 8'h05;
			13'h05bc: data_buf = 8'hcd;
			13'h05bd: data_buf = 8'h4d;
			13'h05be: data_buf = 8'h08;
			13'h05bf: data_buf = 8'h2b;
			13'h05c0: data_buf = 8'h23;
			13'h05c1: data_buf = 8'h7e;
			13'h05c2: data_buf = 8'hfe;
			13'h05c3: data_buf = 8'h61;
			13'h05c4: data_buf = 8'hda;
			13'h05c5: data_buf = 8'hc9;
			13'h05c6: data_buf = 8'h05;
			13'h05c7: data_buf = 8'he6;
			13'h05c8: data_buf = 8'h5f;
			13'h05c9: data_buf = 8'hb9;
			13'h05ca: data_buf = 8'hca;
			13'h05cb: data_buf = 8'haf;
			13'h05cc: data_buf = 8'h05;
			13'h05cd: data_buf = 8'he1;
			13'h05ce: data_buf = 8'hc3;
			13'h05cf: data_buf = 8'h9d;
			13'h05d0: data_buf = 8'h05;
			13'h05d1: data_buf = 8'h48;
			13'h05d2: data_buf = 8'hf1;
			13'h05d3: data_buf = 8'heb;
			13'h05d4: data_buf = 8'hc9;
			13'h05d5: data_buf = 8'heb;
			13'h05d6: data_buf = 8'h79;
			13'h05d7: data_buf = 8'hc1;
			13'h05d8: data_buf = 8'hd1;
			13'h05d9: data_buf = 8'h23;
			13'h05da: data_buf = 8'h12;
			13'h05db: data_buf = 8'h13;
			13'h05dc: data_buf = 8'h0c;
			13'h05dd: data_buf = 8'hd6;
			13'h05de: data_buf = 8'h3a;
			13'h05df: data_buf = 8'hca;
			13'h05e0: data_buf = 8'he7;
			13'h05e1: data_buf = 8'h05;
			13'h05e2: data_buf = 8'hfe;
			13'h05e3: data_buf = 8'h49;
			13'h05e4: data_buf = 8'hc2;
			13'h05e5: data_buf = 8'hea;
			13'h05e6: data_buf = 8'h05;
			13'h05e7: data_buf = 8'h32;
			13'h05e8: data_buf = 8'hf3;
			13'h05e9: data_buf = 8'h80;
			13'h05ea: data_buf = 8'hd6;
			13'h05eb: data_buf = 8'h54;
			13'h05ec: data_buf = 8'hc2;
			13'h05ed: data_buf = 8'h5a;
			13'h05ee: data_buf = 8'h05;
			13'h05ef: data_buf = 8'h47;
			13'h05f0: data_buf = 8'h7e;
			13'h05f1: data_buf = 8'hb7;
			13'h05f2: data_buf = 8'hca;
			13'h05f3: data_buf = 8'h00;
			13'h05f4: data_buf = 8'h06;
			13'h05f5: data_buf = 8'hb8;
			13'h05f6: data_buf = 8'hca;
			13'h05f7: data_buf = 8'hd9;
			13'h05f8: data_buf = 8'h05;
			13'h05f9: data_buf = 8'h23;
			13'h05fa: data_buf = 8'h12;
			13'h05fb: data_buf = 8'h0c;
			13'h05fc: data_buf = 8'h13;
			13'h05fd: data_buf = 8'hc3;
			13'h05fe: data_buf = 8'hf0;
			13'h05ff: data_buf = 8'h05;
			13'h0600: data_buf = 8'h21;
			13'h0601: data_buf = 8'ha5;
			13'h0602: data_buf = 8'h80;
			13'h0603: data_buf = 8'h12;
			13'h0604: data_buf = 8'h13;
			13'h0605: data_buf = 8'h12;
			13'h0606: data_buf = 8'h13;
			13'h0607: data_buf = 8'h12;
			13'h0608: data_buf = 8'hc9;
			13'h0609: data_buf = 8'h3a;
			13'h060a: data_buf = 8'h89;
			13'h060b: data_buf = 8'h80;
			13'h060c: data_buf = 8'hb7;
			13'h060d: data_buf = 8'h3e;
			13'h060e: data_buf = 8'h00;
			13'h060f: data_buf = 8'h32;
			13'h0610: data_buf = 8'h89;
			13'h0611: data_buf = 8'h80;
			13'h0612: data_buf = 8'hc2;
			13'h0613: data_buf = 8'h1d;
			13'h0614: data_buf = 8'h06;
			13'h0615: data_buf = 8'h05;
			13'h0616: data_buf = 8'hca;
			13'h0617: data_buf = 8'h3a;
			13'h0618: data_buf = 8'h06;
			13'h0619: data_buf = 8'hcd;
			13'h061a: data_buf = 8'hce;
			13'h061b: data_buf = 8'h06;
			13'h061c: data_buf = 8'h3e;
			13'h061d: data_buf = 8'h05;
			13'h061e: data_buf = 8'h2b;
			13'h061f: data_buf = 8'hca;
			13'h0620: data_buf = 8'h31;
			13'h0621: data_buf = 8'h06;
			13'h0622: data_buf = 8'h7e;
			13'h0623: data_buf = 8'hcd;
			13'h0624: data_buf = 8'hce;
			13'h0625: data_buf = 8'h06;
			13'h0626: data_buf = 8'hc3;
			13'h0627: data_buf = 8'h43;
			13'h0628: data_buf = 8'h06;
			13'h0629: data_buf = 8'h05;
			13'h062a: data_buf = 8'h2b;
			13'h062b: data_buf = 8'hcd;
			13'h062c: data_buf = 8'hce;
			13'h062d: data_buf = 8'h06;
			13'h062e: data_buf = 8'hc2;
			13'h062f: data_buf = 8'h43;
			13'h0630: data_buf = 8'h06;
			13'h0631: data_buf = 8'hcd;
			13'h0632: data_buf = 8'hce;
			13'h0633: data_buf = 8'h06;
			13'h0634: data_buf = 8'hcd;
			13'h0635: data_buf = 8'hf5;
			13'h0636: data_buf = 8'h0a;
			13'h0637: data_buf = 8'hc3;
			13'h0638: data_buf = 8'h3a;
			13'h0639: data_buf = 8'h06;
			13'h063a: data_buf = 8'h21;
			13'h063b: data_buf = 8'ha6;
			13'h063c: data_buf = 8'h80;
			13'h063d: data_buf = 8'h06;
			13'h063e: data_buf = 8'h01;
			13'h063f: data_buf = 8'haf;
			13'h0640: data_buf = 8'h32;
			13'h0641: data_buf = 8'h89;
			13'h0642: data_buf = 8'h80;
			13'h0643: data_buf = 8'hcd;
			13'h0644: data_buf = 8'hf8;
			13'h0645: data_buf = 8'h06;
			13'h0646: data_buf = 8'h4f;
			13'h0647: data_buf = 8'hfe;
			13'h0648: data_buf = 8'h7f;
			13'h0649: data_buf = 8'hca;
			13'h064a: data_buf = 8'h09;
			13'h064b: data_buf = 8'h06;
			13'h064c: data_buf = 8'h3a;
			13'h064d: data_buf = 8'h89;
			13'h064e: data_buf = 8'h80;
			13'h064f: data_buf = 8'hb7;
			13'h0650: data_buf = 8'hca;
			13'h0651: data_buf = 8'h5c;
			13'h0652: data_buf = 8'h06;
			13'h0653: data_buf = 8'h3e;
			13'h0654: data_buf = 8'h00;
			13'h0655: data_buf = 8'hcd;
			13'h0656: data_buf = 8'hce;
			13'h0657: data_buf = 8'h06;
			13'h0658: data_buf = 8'haf;
			13'h0659: data_buf = 8'h32;
			13'h065a: data_buf = 8'h89;
			13'h065b: data_buf = 8'h80;
			13'h065c: data_buf = 8'h79;
			13'h065d: data_buf = 8'hfe;
			13'h065e: data_buf = 8'h07;
			13'h065f: data_buf = 8'hca;
			13'h0660: data_buf = 8'ha0;
			13'h0661: data_buf = 8'h06;
			13'h0662: data_buf = 8'hfe;
			13'h0663: data_buf = 8'h03;
			13'h0664: data_buf = 8'hcc;
			13'h0665: data_buf = 8'hf5;
			13'h0666: data_buf = 8'h0a;
			13'h0667: data_buf = 8'h37;
			13'h0668: data_buf = 8'hc8;
			13'h0669: data_buf = 8'hfe;
			13'h066a: data_buf = 8'h0d;
			13'h066b: data_buf = 8'hca;
			13'h066c: data_buf = 8'hf0;
			13'h066d: data_buf = 8'h0a;
			13'h066e: data_buf = 8'hfe;
			13'h066f: data_buf = 8'h15;
			13'h0670: data_buf = 8'hca;
			13'h0671: data_buf = 8'h34;
			13'h0672: data_buf = 8'h06;
			13'h0673: data_buf = 8'hfe;
			13'h0674: data_buf = 8'h40;
			13'h0675: data_buf = 8'hca;
			13'h0676: data_buf = 8'h31;
			13'h0677: data_buf = 8'h06;
			13'h0678: data_buf = 8'hfe;
			13'h0679: data_buf = 8'h5f;
			13'h067a: data_buf = 8'hca;
			13'h067b: data_buf = 8'h29;
			13'h067c: data_buf = 8'h06;
			13'h067d: data_buf = 8'hfe;
			13'h067e: data_buf = 8'h08;
			13'h067f: data_buf = 8'hca;
			13'h0680: data_buf = 8'h29;
			13'h0681: data_buf = 8'h06;
			13'h0682: data_buf = 8'hfe;
			13'h0683: data_buf = 8'h12;
			13'h0684: data_buf = 8'hc2;
			13'h0685: data_buf = 8'h9b;
			13'h0686: data_buf = 8'h06;
			13'h0687: data_buf = 8'hc5;
			13'h0688: data_buf = 8'hd5;
			13'h0689: data_buf = 8'he5;
			13'h068a: data_buf = 8'h36;
			13'h068b: data_buf = 8'h00;
			13'h068c: data_buf = 8'hcd;
			13'h068d: data_buf = 8'h9f;
			13'h068e: data_buf = 8'h1c;
			13'h068f: data_buf = 8'h21;
			13'h0690: data_buf = 8'ha6;
			13'h0691: data_buf = 8'h80;
			13'h0692: data_buf = 8'hcd;
			13'h0693: data_buf = 8'h93;
			13'h0694: data_buf = 8'h11;
			13'h0695: data_buf = 8'he1;
			13'h0696: data_buf = 8'hd1;
			13'h0697: data_buf = 8'hc1;
			13'h0698: data_buf = 8'hc3;
			13'h0699: data_buf = 8'h43;
			13'h069a: data_buf = 8'h06;
			13'h069b: data_buf = 8'hfe;
			13'h069c: data_buf = 8'h20;
			13'h069d: data_buf = 8'hda;
			13'h069e: data_buf = 8'h43;
			13'h069f: data_buf = 8'h06;
			13'h06a0: data_buf = 8'h78;
			13'h06a1: data_buf = 8'hfe;
			13'h06a2: data_buf = 8'h49;
			13'h06a3: data_buf = 8'h3e;
			13'h06a4: data_buf = 8'h07;
			13'h06a5: data_buf = 8'hd2;
			13'h06a6: data_buf = 8'hb5;
			13'h06a7: data_buf = 8'h06;
			13'h06a8: data_buf = 8'h79;
			13'h06a9: data_buf = 8'h71;
			13'h06aa: data_buf = 8'h32;
			13'h06ab: data_buf = 8'h11;
			13'h06ac: data_buf = 8'h81;
			13'h06ad: data_buf = 8'h23;
			13'h06ae: data_buf = 8'h04;
			13'h06af: data_buf = 8'hcd;
			13'h06b0: data_buf = 8'hce;
			13'h06b1: data_buf = 8'h06;
			13'h06b2: data_buf = 8'hc3;
			13'h06b3: data_buf = 8'h43;
			13'h06b4: data_buf = 8'h06;
			13'h06b5: data_buf = 8'hcd;
			13'h06b6: data_buf = 8'hce;
			13'h06b7: data_buf = 8'h06;
			13'h06b8: data_buf = 8'h3e;
			13'h06b9: data_buf = 8'h08;
			13'h06ba: data_buf = 8'hc3;
			13'h06bb: data_buf = 8'haf;
			13'h06bc: data_buf = 8'h06;
			13'h06bd: data_buf = 8'h7c;
			13'h06be: data_buf = 8'h92;
			13'h06bf: data_buf = 8'hc0;
			13'h06c0: data_buf = 8'h7d;
			13'h06c1: data_buf = 8'h93;
			13'h06c2: data_buf = 8'hc9;
			13'h06c3: data_buf = 8'h7e;
			13'h06c4: data_buf = 8'he3;
			13'h06c5: data_buf = 8'hbe;
			13'h06c6: data_buf = 8'h23;
			13'h06c7: data_buf = 8'he3;
			13'h06c8: data_buf = 8'hca;
			13'h06c9: data_buf = 8'h4d;
			13'h06ca: data_buf = 8'h08;
			13'h06cb: data_buf = 8'hc3;
			13'h06cc: data_buf = 8'hf5;
			13'h06cd: data_buf = 8'h03;
			13'h06ce: data_buf = 8'hf5;
			13'h06cf: data_buf = 8'h3a;
			13'h06d0: data_buf = 8'h8a;
			13'h06d1: data_buf = 8'h80;
			13'h06d2: data_buf = 8'hb7;
			13'h06d3: data_buf = 8'hc2;
			13'h06d4: data_buf = 8'hc8;
			13'h06d5: data_buf = 8'h11;
			13'h06d6: data_buf = 8'hf1;
			13'h06d7: data_buf = 8'hc5;
			13'h06d8: data_buf = 8'hf5;
			13'h06d9: data_buf = 8'hfe;
			13'h06da: data_buf = 8'h20;
			13'h06db: data_buf = 8'hda;
			13'h06dc: data_buf = 8'hf2;
			13'h06dd: data_buf = 8'h06;
			13'h06de: data_buf = 8'h3a;
			13'h06df: data_buf = 8'h87;
			13'h06e0: data_buf = 8'h80;
			13'h06e1: data_buf = 8'h47;
			13'h06e2: data_buf = 8'h3a;
			13'h06e3: data_buf = 8'hf0;
			13'h06e4: data_buf = 8'h80;
			13'h06e5: data_buf = 8'h04;
			13'h06e6: data_buf = 8'hca;
			13'h06e7: data_buf = 8'hee;
			13'h06e8: data_buf = 8'h06;
			13'h06e9: data_buf = 8'h05;
			13'h06ea: data_buf = 8'hb8;
			13'h06eb: data_buf = 8'hcc;
			13'h06ec: data_buf = 8'hf5;
			13'h06ed: data_buf = 8'h0a;
			13'h06ee: data_buf = 8'h3c;
			13'h06ef: data_buf = 8'h32;
			13'h06f0: data_buf = 8'hf0;
			13'h06f1: data_buf = 8'h80;
			13'h06f2: data_buf = 8'hf1;
			13'h06f3: data_buf = 8'hc1;
			13'h06f4: data_buf = 8'hcd;
			13'h06f5: data_buf = 8'h8a;
			13'h06f6: data_buf = 8'h1c;
			13'h06f7: data_buf = 8'hc9;
			13'h06f8: data_buf = 8'hcd;
			13'h06f9: data_buf = 8'h52;
			13'h06fa: data_buf = 8'h1b;
			13'h06fb: data_buf = 8'he6;
			13'h06fc: data_buf = 8'h7f;
			13'h06fd: data_buf = 8'hfe;
			13'h06fe: data_buf = 8'h0f;
			13'h06ff: data_buf = 8'hc0;
			13'h0700: data_buf = 8'h3a;
			13'h0701: data_buf = 8'h8a;
			13'h0702: data_buf = 8'h80;
			13'h0703: data_buf = 8'h2f;
			13'h0704: data_buf = 8'h32;
			13'h0705: data_buf = 8'h8a;
			13'h0706: data_buf = 8'h80;
			13'h0707: data_buf = 8'haf;
			13'h0708: data_buf = 8'hc9;
			13'h0709: data_buf = 8'hcd;
			13'h070a: data_buf = 8'h19;
			13'h070b: data_buf = 8'h09;
			13'h070c: data_buf = 8'hc0;
			13'h070d: data_buf = 8'hc1;
			13'h070e: data_buf = 8'hcd;
			13'h070f: data_buf = 8'he1;
			13'h0710: data_buf = 8'h04;
			13'h0711: data_buf = 8'hc5;
			13'h0712: data_buf = 8'hcd;
			13'h0713: data_buf = 8'h5f;
			13'h0714: data_buf = 8'h07;
			13'h0715: data_buf = 8'he1;
			13'h0716: data_buf = 8'h4e;
			13'h0717: data_buf = 8'h23;
			13'h0718: data_buf = 8'h46;
			13'h0719: data_buf = 8'h23;
			13'h071a: data_buf = 8'h78;
			13'h071b: data_buf = 8'hb1;
			13'h071c: data_buf = 8'hca;
			13'h071d: data_buf = 8'h40;
			13'h071e: data_buf = 8'h04;
			13'h071f: data_buf = 8'hcd;
			13'h0720: data_buf = 8'h68;
			13'h0721: data_buf = 8'h07;
			13'h0722: data_buf = 8'hcd;
			13'h0723: data_buf = 8'h78;
			13'h0724: data_buf = 8'h08;
			13'h0725: data_buf = 8'hc5;
			13'h0726: data_buf = 8'hcd;
			13'h0727: data_buf = 8'hf5;
			13'h0728: data_buf = 8'h0a;
			13'h0729: data_buf = 8'h5e;
			13'h072a: data_buf = 8'h23;
			13'h072b: data_buf = 8'h56;
			13'h072c: data_buf = 8'h23;
			13'h072d: data_buf = 8'he5;
			13'h072e: data_buf = 8'heb;
			13'h072f: data_buf = 8'hcd;
			13'h0730: data_buf = 8'h36;
			13'h0731: data_buf = 8'h18;
			13'h0732: data_buf = 8'h3e;
			13'h0733: data_buf = 8'h20;
			13'h0734: data_buf = 8'he1;
			13'h0735: data_buf = 8'hcd;
			13'h0736: data_buf = 8'hce;
			13'h0737: data_buf = 8'h06;
			13'h0738: data_buf = 8'h7e;
			13'h0739: data_buf = 8'hb7;
			13'h073a: data_buf = 8'h23;
			13'h073b: data_buf = 8'hca;
			13'h073c: data_buf = 8'h15;
			13'h073d: data_buf = 8'h07;
			13'h073e: data_buf = 8'hf2;
			13'h073f: data_buf = 8'h35;
			13'h0740: data_buf = 8'h07;
			13'h0741: data_buf = 8'hd6;
			13'h0742: data_buf = 8'h7f;
			13'h0743: data_buf = 8'h4f;
			13'h0744: data_buf = 8'h11;
			13'h0745: data_buf = 8'h7e;
			13'h0746: data_buf = 8'h01;
			13'h0747: data_buf = 8'h1a;
			13'h0748: data_buf = 8'h13;
			13'h0749: data_buf = 8'hb7;
			13'h074a: data_buf = 8'hf2;
			13'h074b: data_buf = 8'h47;
			13'h074c: data_buf = 8'h07;
			13'h074d: data_buf = 8'h0d;
			13'h074e: data_buf = 8'hc2;
			13'h074f: data_buf = 8'h47;
			13'h0750: data_buf = 8'h07;
			13'h0751: data_buf = 8'he6;
			13'h0752: data_buf = 8'h7f;
			13'h0753: data_buf = 8'hcd;
			13'h0754: data_buf = 8'hce;
			13'h0755: data_buf = 8'h06;
			13'h0756: data_buf = 8'h1a;
			13'h0757: data_buf = 8'h13;
			13'h0758: data_buf = 8'hb7;
			13'h0759: data_buf = 8'hf2;
			13'h075a: data_buf = 8'h51;
			13'h075b: data_buf = 8'h07;
			13'h075c: data_buf = 8'hc3;
			13'h075d: data_buf = 8'h38;
			13'h075e: data_buf = 8'h07;
			13'h075f: data_buf = 8'he5;
			13'h0760: data_buf = 8'h2a;
			13'h0761: data_buf = 8'h8d;
			13'h0762: data_buf = 8'h80;
			13'h0763: data_buf = 8'h22;
			13'h0764: data_buf = 8'h8b;
			13'h0765: data_buf = 8'h80;
			13'h0766: data_buf = 8'he1;
			13'h0767: data_buf = 8'hc9;
			13'h0768: data_buf = 8'he5;
			13'h0769: data_buf = 8'hd5;
			13'h076a: data_buf = 8'h2a;
			13'h076b: data_buf = 8'h8b;
			13'h076c: data_buf = 8'h80;
			13'h076d: data_buf = 8'h11;
			13'h076e: data_buf = 8'hff;
			13'h076f: data_buf = 8'hff;
			13'h0770: data_buf = 8'hed;
			13'h0771: data_buf = 8'h5a;
			13'h0772: data_buf = 8'h22;
			13'h0773: data_buf = 8'h8b;
			13'h0774: data_buf = 8'h80;
			13'h0775: data_buf = 8'hd1;
			13'h0776: data_buf = 8'he1;
			13'h0777: data_buf = 8'hf0;
			13'h0778: data_buf = 8'he5;
			13'h0779: data_buf = 8'h2a;
			13'h077a: data_buf = 8'h8d;
			13'h077b: data_buf = 8'h80;
			13'h077c: data_buf = 8'h22;
			13'h077d: data_buf = 8'h8b;
			13'h077e: data_buf = 8'h80;
			13'h077f: data_buf = 8'hcd;
			13'h0780: data_buf = 8'h52;
			13'h0781: data_buf = 8'h1b;
			13'h0782: data_buf = 8'hfe;
			13'h0783: data_buf = 8'h03;
			13'h0784: data_buf = 8'hca;
			13'h0785: data_buf = 8'h8b;
			13'h0786: data_buf = 8'h07;
			13'h0787: data_buf = 8'he1;
			13'h0788: data_buf = 8'hc3;
			13'h0789: data_buf = 8'h68;
			13'h078a: data_buf = 8'h07;
			13'h078b: data_buf = 8'h2a;
			13'h078c: data_buf = 8'h8d;
			13'h078d: data_buf = 8'h80;
			13'h078e: data_buf = 8'h22;
			13'h078f: data_buf = 8'h8b;
			13'h0790: data_buf = 8'h80;
			13'h0791: data_buf = 8'hc3;
			13'h0792: data_buf = 8'hbf;
			13'h0793: data_buf = 8'h00;
			13'h0794: data_buf = 8'h3e;
			13'h0795: data_buf = 8'h64;
			13'h0796: data_buf = 8'h32;
			13'h0797: data_buf = 8'h10;
			13'h0798: data_buf = 8'h81;
			13'h0799: data_buf = 8'hcd;
			13'h079a: data_buf = 8'hfb;
			13'h079b: data_buf = 8'h09;
			13'h079c: data_buf = 8'hc1;
			13'h079d: data_buf = 8'he5;
			13'h079e: data_buf = 8'hcd;
			13'h079f: data_buf = 8'he4;
			13'h07a0: data_buf = 8'h09;
			13'h07a1: data_buf = 8'h22;
			13'h07a2: data_buf = 8'h0c;
			13'h07a3: data_buf = 8'h81;
			13'h07a4: data_buf = 8'h21;
			13'h07a5: data_buf = 8'h02;
			13'h07a6: data_buf = 8'h00;
			13'h07a7: data_buf = 8'h39;
			13'h07a8: data_buf = 8'hcd;
			13'h07a9: data_buf = 8'ha2;
			13'h07aa: data_buf = 8'h03;
			13'h07ab: data_buf = 8'hd1;
			13'h07ac: data_buf = 8'hc2;
			13'h07ad: data_buf = 8'hc4;
			13'h07ae: data_buf = 8'h07;
			13'h07af: data_buf = 8'h09;
			13'h07b0: data_buf = 8'hd5;
			13'h07b1: data_buf = 8'h2b;
			13'h07b2: data_buf = 8'h56;
			13'h07b3: data_buf = 8'h2b;
			13'h07b4: data_buf = 8'h5e;
			13'h07b5: data_buf = 8'h23;
			13'h07b6: data_buf = 8'h23;
			13'h07b7: data_buf = 8'he5;
			13'h07b8: data_buf = 8'h2a;
			13'h07b9: data_buf = 8'h0c;
			13'h07ba: data_buf = 8'h81;
			13'h07bb: data_buf = 8'hcd;
			13'h07bc: data_buf = 8'hbd;
			13'h07bd: data_buf = 8'h06;
			13'h07be: data_buf = 8'he1;
			13'h07bf: data_buf = 8'hc2;
			13'h07c0: data_buf = 8'ha8;
			13'h07c1: data_buf = 8'h07;
			13'h07c2: data_buf = 8'hd1;
			13'h07c3: data_buf = 8'hf9;
			13'h07c4: data_buf = 8'heb;
			13'h07c5: data_buf = 8'h0e;
			13'h07c6: data_buf = 8'h08;
			13'h07c7: data_buf = 8'hcd;
			13'h07c8: data_buf = 8'hd2;
			13'h07c9: data_buf = 8'h03;
			13'h07ca: data_buf = 8'he5;
			13'h07cb: data_buf = 8'h2a;
			13'h07cc: data_buf = 8'h0c;
			13'h07cd: data_buf = 8'h81;
			13'h07ce: data_buf = 8'he3;
			13'h07cf: data_buf = 8'he5;
			13'h07d0: data_buf = 8'h2a;
			13'h07d1: data_buf = 8'ha1;
			13'h07d2: data_buf = 8'h80;
			13'h07d3: data_buf = 8'he3;
			13'h07d4: data_buf = 8'hcd;
			13'h07d5: data_buf = 8'hbd;
			13'h07d6: data_buf = 8'h0c;
			13'h07d7: data_buf = 8'hcd;
			13'h07d8: data_buf = 8'hc3;
			13'h07d9: data_buf = 8'h06;
			13'h07da: data_buf = 8'ha6;
			13'h07db: data_buf = 8'hcd;
			13'h07dc: data_buf = 8'hba;
			13'h07dd: data_buf = 8'h0c;
			13'h07de: data_buf = 8'he5;
			13'h07df: data_buf = 8'hcd;
			13'h07e0: data_buf = 8'he8;
			13'h07e1: data_buf = 8'h16;
			13'h07e2: data_buf = 8'he1;
			13'h07e3: data_buf = 8'hc5;
			13'h07e4: data_buf = 8'hd5;
			13'h07e5: data_buf = 8'h01;
			13'h07e6: data_buf = 8'h00;
			13'h07e7: data_buf = 8'h81;
			13'h07e8: data_buf = 8'h51;
			13'h07e9: data_buf = 8'h5a;
			13'h07ea: data_buf = 8'h7e;
			13'h07eb: data_buf = 8'hfe;
			13'h07ec: data_buf = 8'hab;
			13'h07ed: data_buf = 8'h3e;
			13'h07ee: data_buf = 8'h01;
			13'h07ef: data_buf = 8'hc2;
			13'h07f0: data_buf = 8'h00;
			13'h07f1: data_buf = 8'h08;
			13'h07f2: data_buf = 8'hcd;
			13'h07f3: data_buf = 8'h4d;
			13'h07f4: data_buf = 8'h08;
			13'h07f5: data_buf = 8'hcd;
			13'h07f6: data_buf = 8'hba;
			13'h07f7: data_buf = 8'h0c;
			13'h07f8: data_buf = 8'he5;
			13'h07f9: data_buf = 8'hcd;
			13'h07fa: data_buf = 8'he8;
			13'h07fb: data_buf = 8'h16;
			13'h07fc: data_buf = 8'hcd;
			13'h07fd: data_buf = 8'h9c;
			13'h07fe: data_buf = 8'h16;
			13'h07ff: data_buf = 8'he1;
			13'h0800: data_buf = 8'hc5;
			13'h0801: data_buf = 8'hd5;
			13'h0802: data_buf = 8'hf5;
			13'h0803: data_buf = 8'h33;
			13'h0804: data_buf = 8'he5;
			13'h0805: data_buf = 8'h2a;
			13'h0806: data_buf = 8'h13;
			13'h0807: data_buf = 8'h81;
			13'h0808: data_buf = 8'he3;
			13'h0809: data_buf = 8'h06;
			13'h080a: data_buf = 8'h81;
			13'h080b: data_buf = 8'hc5;
			13'h080c: data_buf = 8'h33;
			13'h080d: data_buf = 8'hcd;
			13'h080e: data_buf = 8'h78;
			13'h080f: data_buf = 8'h08;
			13'h0810: data_buf = 8'h22;
			13'h0811: data_buf = 8'h13;
			13'h0812: data_buf = 8'h81;
			13'h0813: data_buf = 8'h7e;
			13'h0814: data_buf = 8'hfe;
			13'h0815: data_buf = 8'h3a;
			13'h0816: data_buf = 8'hca;
			13'h0817: data_buf = 8'h2d;
			13'h0818: data_buf = 8'h08;
			13'h0819: data_buf = 8'hb7;
			13'h081a: data_buf = 8'hc2;
			13'h081b: data_buf = 8'hf5;
			13'h081c: data_buf = 8'h03;
			13'h081d: data_buf = 8'h23;
			13'h081e: data_buf = 8'h7e;
			13'h081f: data_buf = 8'h23;
			13'h0820: data_buf = 8'hb6;
			13'h0821: data_buf = 8'hca;
			13'h0822: data_buf = 8'h9f;
			13'h0823: data_buf = 8'h08;
			13'h0824: data_buf = 8'h23;
			13'h0825: data_buf = 8'h5e;
			13'h0826: data_buf = 8'h23;
			13'h0827: data_buf = 8'h56;
			13'h0828: data_buf = 8'heb;
			13'h0829: data_buf = 8'h22;
			13'h082a: data_buf = 8'ha1;
			13'h082b: data_buf = 8'h80;
			13'h082c: data_buf = 8'heb;
			13'h082d: data_buf = 8'hcd;
			13'h082e: data_buf = 8'h4d;
			13'h082f: data_buf = 8'h08;
			13'h0830: data_buf = 8'h11;
			13'h0831: data_buf = 8'h0d;
			13'h0832: data_buf = 8'h08;
			13'h0833: data_buf = 8'hd5;
			13'h0834: data_buf = 8'hc8;
			13'h0835: data_buf = 8'hd6;
			13'h0836: data_buf = 8'h80;
			13'h0837: data_buf = 8'hda;
			13'h0838: data_buf = 8'hfb;
			13'h0839: data_buf = 8'h09;
			13'h083a: data_buf = 8'hfe;
			13'h083b: data_buf = 8'h25;
			13'h083c: data_buf = 8'hd2;
			13'h083d: data_buf = 8'hf5;
			13'h083e: data_buf = 8'h03;
			13'h083f: data_buf = 8'h07;
			13'h0840: data_buf = 8'h4f;
			13'h0841: data_buf = 8'h06;
			13'h0842: data_buf = 8'h00;
			13'h0843: data_buf = 8'heb;
			13'h0844: data_buf = 8'h21;
			13'h0845: data_buf = 8'h9d;
			13'h0846: data_buf = 8'h02;
			13'h0847: data_buf = 8'h09;
			13'h0848: data_buf = 8'h4e;
			13'h0849: data_buf = 8'h23;
			13'h084a: data_buf = 8'h46;
			13'h084b: data_buf = 8'hc5;
			13'h084c: data_buf = 8'heb;
			13'h084d: data_buf = 8'h23;
			13'h084e: data_buf = 8'h7e;
			13'h084f: data_buf = 8'hfe;
			13'h0850: data_buf = 8'h3a;
			13'h0851: data_buf = 8'hd0;
			13'h0852: data_buf = 8'hfe;
			13'h0853: data_buf = 8'h20;
			13'h0854: data_buf = 8'hca;
			13'h0855: data_buf = 8'h4d;
			13'h0856: data_buf = 8'h08;
			13'h0857: data_buf = 8'hfe;
			13'h0858: data_buf = 8'h30;
			13'h0859: data_buf = 8'h3f;
			13'h085a: data_buf = 8'h3c;
			13'h085b: data_buf = 8'h3d;
			13'h085c: data_buf = 8'hc9;
			13'h085d: data_buf = 8'heb;
			13'h085e: data_buf = 8'h2a;
			13'h085f: data_buf = 8'ha3;
			13'h0860: data_buf = 8'h80;
			13'h0861: data_buf = 8'hca;
			13'h0862: data_buf = 8'h72;
			13'h0863: data_buf = 8'h08;
			13'h0864: data_buf = 8'heb;
			13'h0865: data_buf = 8'hcd;
			13'h0866: data_buf = 8'h19;
			13'h0867: data_buf = 8'h09;
			13'h0868: data_buf = 8'he5;
			13'h0869: data_buf = 8'hcd;
			13'h086a: data_buf = 8'he1;
			13'h086b: data_buf = 8'h04;
			13'h086c: data_buf = 8'h60;
			13'h086d: data_buf = 8'h69;
			13'h086e: data_buf = 8'hd1;
			13'h086f: data_buf = 8'hd2;
			13'h0870: data_buf = 8'hba;
			13'h0871: data_buf = 8'h09;
			13'h0872: data_buf = 8'h2b;
			13'h0873: data_buf = 8'h22;
			13'h0874: data_buf = 8'h21;
			13'h0875: data_buf = 8'h81;
			13'h0876: data_buf = 8'heb;
			13'h0877: data_buf = 8'hc9;
			13'h0878: data_buf = 8'hdf;
			13'h0879: data_buf = 8'hc8;
			13'h087a: data_buf = 8'hd7;
			13'h087b: data_buf = 8'hfe;
			13'h087c: data_buf = 8'h1b;
			13'h087d: data_buf = 8'h28;
			13'h087e: data_buf = 8'h11;
			13'h087f: data_buf = 8'hfe;
			13'h0880: data_buf = 8'h03;
			13'h0881: data_buf = 8'h28;
			13'h0882: data_buf = 8'h0d;
			13'h0883: data_buf = 8'hfe;
			13'h0884: data_buf = 8'h13;
			13'h0885: data_buf = 8'hc0;
			13'h0886: data_buf = 8'hd7;
			13'h0887: data_buf = 8'hfe;
			13'h0888: data_buf = 8'h11;
			13'h0889: data_buf = 8'hc8;
			13'h088a: data_buf = 8'hfe;
			13'h088b: data_buf = 8'h03;
			13'h088c: data_buf = 8'h28;
			13'h088d: data_buf = 8'h07;
			13'h088e: data_buf = 8'h18;
			13'h088f: data_buf = 8'hf6;
			13'h0890: data_buf = 8'h3e;
			13'h0891: data_buf = 8'hff;
			13'h0892: data_buf = 8'h32;
			13'h0893: data_buf = 8'h92;
			13'h0894: data_buf = 8'h80;
			13'h0895: data_buf = 8'hc0;
			13'h0896: data_buf = 8'hf6;
			13'h0897: data_buf = 8'hc0;
			13'h0898: data_buf = 8'h22;
			13'h0899: data_buf = 8'h13;
			13'h089a: data_buf = 8'h81;
			13'h089b: data_buf = 8'h21;
			13'h089c: data_buf = 8'hf6;
			13'h089d: data_buf = 8'hff;
			13'h089e: data_buf = 8'hc1;
			13'h089f: data_buf = 8'h2a;
			13'h08a0: data_buf = 8'ha1;
			13'h08a1: data_buf = 8'h80;
			13'h08a2: data_buf = 8'hf5;
			13'h08a3: data_buf = 8'h7d;
			13'h08a4: data_buf = 8'ha4;
			13'h08a5: data_buf = 8'h3c;
			13'h08a6: data_buf = 8'hca;
			13'h08a7: data_buf = 8'hb2;
			13'h08a8: data_buf = 8'h08;
			13'h08a9: data_buf = 8'h22;
			13'h08aa: data_buf = 8'h17;
			13'h08ab: data_buf = 8'h81;
			13'h08ac: data_buf = 8'h2a;
			13'h08ad: data_buf = 8'h13;
			13'h08ae: data_buf = 8'h81;
			13'h08af: data_buf = 8'h22;
			13'h08b0: data_buf = 8'h19;
			13'h08b1: data_buf = 8'h81;
			13'h08b2: data_buf = 8'haf;
			13'h08b3: data_buf = 8'h32;
			13'h08b4: data_buf = 8'h8a;
			13'h08b5: data_buf = 8'h80;
			13'h08b6: data_buf = 8'hcd;
			13'h08b7: data_buf = 8'he8;
			13'h08b8: data_buf = 8'h0a;
			13'h08b9: data_buf = 8'hf1;
			13'h08ba: data_buf = 8'h21;
			13'h08bb: data_buf = 8'h98;
			13'h08bc: data_buf = 8'h03;
			13'h08bd: data_buf = 8'hc2;
			13'h08be: data_buf = 8'h29;
			13'h08bf: data_buf = 8'h04;
			13'h08c0: data_buf = 8'hc3;
			13'h08c1: data_buf = 8'h40;
			13'h08c2: data_buf = 8'h04;
			13'h08c3: data_buf = 8'h2a;
			13'h08c4: data_buf = 8'h19;
			13'h08c5: data_buf = 8'h81;
			13'h08c6: data_buf = 8'h7c;
			13'h08c7: data_buf = 8'hb5;
			13'h08c8: data_buf = 8'h1e;
			13'h08c9: data_buf = 8'h20;
			13'h08ca: data_buf = 8'hca;
			13'h08cb: data_buf = 8'h09;
			13'h08cc: data_buf = 8'h04;
			13'h08cd: data_buf = 8'heb;
			13'h08ce: data_buf = 8'h2a;
			13'h08cf: data_buf = 8'h17;
			13'h08d0: data_buf = 8'h81;
			13'h08d1: data_buf = 8'h22;
			13'h08d2: data_buf = 8'ha1;
			13'h08d3: data_buf = 8'h80;
			13'h08d4: data_buf = 8'heb;
			13'h08d5: data_buf = 8'hc9;
			13'h08d6: data_buf = 8'hcd;
			13'h08d7: data_buf = 8'h1b;
			13'h08d8: data_buf = 8'h14;
			13'h08d9: data_buf = 8'hc0;
			13'h08da: data_buf = 8'h32;
			13'h08db: data_buf = 8'h86;
			13'h08dc: data_buf = 8'h80;
			13'h08dd: data_buf = 8'hc9;
			13'h08de: data_buf = 8'he5;
			13'h08df: data_buf = 8'h2a;
			13'h08e0: data_buf = 8'h8f;
			13'h08e1: data_buf = 8'h80;
			13'h08e2: data_buf = 8'h06;
			13'h08e3: data_buf = 8'h00;
			13'h08e4: data_buf = 8'h4f;
			13'h08e5: data_buf = 8'h09;
			13'h08e6: data_buf = 8'h22;
			13'h08e7: data_buf = 8'h8f;
			13'h08e8: data_buf = 8'h80;
			13'h08e9: data_buf = 8'he1;
			13'h08ea: data_buf = 8'hc9;
			13'h08eb: data_buf = 8'h7e;
			13'h08ec: data_buf = 8'hfe;
			13'h08ed: data_buf = 8'h41;
			13'h08ee: data_buf = 8'hd8;
			13'h08ef: data_buf = 8'hfe;
			13'h08f0: data_buf = 8'h5b;
			13'h08f1: data_buf = 8'h3f;
			13'h08f2: data_buf = 8'hc9;
			13'h08f3: data_buf = 8'hcd;
			13'h08f4: data_buf = 8'h4d;
			13'h08f5: data_buf = 8'h08;
			13'h08f6: data_buf = 8'hcd;
			13'h08f7: data_buf = 8'hba;
			13'h08f8: data_buf = 8'h0c;
			13'h08f9: data_buf = 8'hcd;
			13'h08fa: data_buf = 8'h9c;
			13'h08fb: data_buf = 8'h16;
			13'h08fc: data_buf = 8'hfa;
			13'h08fd: data_buf = 8'h14;
			13'h08fe: data_buf = 8'h09;
			13'h08ff: data_buf = 8'h3a;
			13'h0900: data_buf = 8'h2c;
			13'h0901: data_buf = 8'h81;
			13'h0902: data_buf = 8'hfe;
			13'h0903: data_buf = 8'h90;
			13'h0904: data_buf = 8'hda;
			13'h0905: data_buf = 8'h44;
			13'h0906: data_buf = 8'h17;
			13'h0907: data_buf = 8'h01;
			13'h0908: data_buf = 8'h80;
			13'h0909: data_buf = 8'h90;
			13'h090a: data_buf = 8'h11;
			13'h090b: data_buf = 8'h00;
			13'h090c: data_buf = 8'h00;
			13'h090d: data_buf = 8'he5;
			13'h090e: data_buf = 8'hcd;
			13'h090f: data_buf = 8'h17;
			13'h0910: data_buf = 8'h17;
			13'h0911: data_buf = 8'he1;
			13'h0912: data_buf = 8'h51;
			13'h0913: data_buf = 8'hc8;
			13'h0914: data_buf = 8'h1e;
			13'h0915: data_buf = 8'h08;
			13'h0916: data_buf = 8'hc3;
			13'h0917: data_buf = 8'h09;
			13'h0918: data_buf = 8'h04;
			13'h0919: data_buf = 8'h2b;
			13'h091a: data_buf = 8'h11;
			13'h091b: data_buf = 8'h00;
			13'h091c: data_buf = 8'h00;
			13'h091d: data_buf = 8'hcd;
			13'h091e: data_buf = 8'h4d;
			13'h091f: data_buf = 8'h08;
			13'h0920: data_buf = 8'hd0;
			13'h0921: data_buf = 8'he5;
			13'h0922: data_buf = 8'hf5;
			13'h0923: data_buf = 8'h21;
			13'h0924: data_buf = 8'h98;
			13'h0925: data_buf = 8'h19;
			13'h0926: data_buf = 8'hcd;
			13'h0927: data_buf = 8'hbd;
			13'h0928: data_buf = 8'h06;
			13'h0929: data_buf = 8'hda;
			13'h092a: data_buf = 8'hf5;
			13'h092b: data_buf = 8'h03;
			13'h092c: data_buf = 8'h62;
			13'h092d: data_buf = 8'h6b;
			13'h092e: data_buf = 8'h19;
			13'h092f: data_buf = 8'h29;
			13'h0930: data_buf = 8'h19;
			13'h0931: data_buf = 8'h29;
			13'h0932: data_buf = 8'hf1;
			13'h0933: data_buf = 8'hd6;
			13'h0934: data_buf = 8'h30;
			13'h0935: data_buf = 8'h5f;
			13'h0936: data_buf = 8'h16;
			13'h0937: data_buf = 8'h00;
			13'h0938: data_buf = 8'h19;
			13'h0939: data_buf = 8'heb;
			13'h093a: data_buf = 8'he1;
			13'h093b: data_buf = 8'hc3;
			13'h093c: data_buf = 8'h1d;
			13'h093d: data_buf = 8'h09;
			13'h093e: data_buf = 8'hca;
			13'h093f: data_buf = 8'h11;
			13'h0940: data_buf = 8'h05;
			13'h0941: data_buf = 8'hcd;
			13'h0942: data_buf = 8'hf6;
			13'h0943: data_buf = 8'h08;
			13'h0944: data_buf = 8'h2b;
			13'h0945: data_buf = 8'hcd;
			13'h0946: data_buf = 8'h4d;
			13'h0947: data_buf = 8'h08;
			13'h0948: data_buf = 8'he5;
			13'h0949: data_buf = 8'h2a;
			13'h094a: data_buf = 8'hf4;
			13'h094b: data_buf = 8'h80;
			13'h094c: data_buf = 8'hca;
			13'h094d: data_buf = 8'h61;
			13'h094e: data_buf = 8'h09;
			13'h094f: data_buf = 8'he1;
			13'h0950: data_buf = 8'hcd;
			13'h0951: data_buf = 8'hc3;
			13'h0952: data_buf = 8'h06;
			13'h0953: data_buf = 8'h2c;
			13'h0954: data_buf = 8'hd5;
			13'h0955: data_buf = 8'hcd;
			13'h0956: data_buf = 8'hf6;
			13'h0957: data_buf = 8'h08;
			13'h0958: data_buf = 8'h2b;
			13'h0959: data_buf = 8'hcd;
			13'h095a: data_buf = 8'h4d;
			13'h095b: data_buf = 8'h08;
			13'h095c: data_buf = 8'hc2;
			13'h095d: data_buf = 8'hf5;
			13'h095e: data_buf = 8'h03;
			13'h095f: data_buf = 8'he3;
			13'h0960: data_buf = 8'heb;
			13'h0961: data_buf = 8'h7d;
			13'h0962: data_buf = 8'h93;
			13'h0963: data_buf = 8'h5f;
			13'h0964: data_buf = 8'h7c;
			13'h0965: data_buf = 8'h9a;
			13'h0966: data_buf = 8'h57;
			13'h0967: data_buf = 8'hda;
			13'h0968: data_buf = 8'hea;
			13'h0969: data_buf = 8'h03;
			13'h096a: data_buf = 8'he5;
			13'h096b: data_buf = 8'h2a;
			13'h096c: data_buf = 8'h1b;
			13'h096d: data_buf = 8'h81;
			13'h096e: data_buf = 8'h01;
			13'h096f: data_buf = 8'h28;
			13'h0970: data_buf = 8'h00;
			13'h0971: data_buf = 8'h09;
			13'h0972: data_buf = 8'hcd;
			13'h0973: data_buf = 8'hbd;
			13'h0974: data_buf = 8'h06;
			13'h0975: data_buf = 8'hd2;
			13'h0976: data_buf = 8'hea;
			13'h0977: data_buf = 8'h03;
			13'h0978: data_buf = 8'heb;
			13'h0979: data_buf = 8'h22;
			13'h097a: data_buf = 8'h9f;
			13'h097b: data_buf = 8'h80;
			13'h097c: data_buf = 8'he1;
			13'h097d: data_buf = 8'h22;
			13'h097e: data_buf = 8'hf4;
			13'h097f: data_buf = 8'h80;
			13'h0980: data_buf = 8'he1;
			13'h0981: data_buf = 8'hc3;
			13'h0982: data_buf = 8'h11;
			13'h0983: data_buf = 8'h05;
			13'h0984: data_buf = 8'hca;
			13'h0985: data_buf = 8'h0d;
			13'h0986: data_buf = 8'h05;
			13'h0987: data_buf = 8'hcd;
			13'h0988: data_buf = 8'h11;
			13'h0989: data_buf = 8'h05;
			13'h098a: data_buf = 8'h01;
			13'h098b: data_buf = 8'h0d;
			13'h098c: data_buf = 8'h08;
			13'h098d: data_buf = 8'hc3;
			13'h098e: data_buf = 8'ha0;
			13'h098f: data_buf = 8'h09;
			13'h0990: data_buf = 8'h0e;
			13'h0991: data_buf = 8'h03;
			13'h0992: data_buf = 8'hcd;
			13'h0993: data_buf = 8'hd2;
			13'h0994: data_buf = 8'h03;
			13'h0995: data_buf = 8'hc1;
			13'h0996: data_buf = 8'he5;
			13'h0997: data_buf = 8'he5;
			13'h0998: data_buf = 8'h2a;
			13'h0999: data_buf = 8'ha1;
			13'h099a: data_buf = 8'h80;
			13'h099b: data_buf = 8'he3;
			13'h099c: data_buf = 8'h3e;
			13'h099d: data_buf = 8'h8c;
			13'h099e: data_buf = 8'hf5;
			13'h099f: data_buf = 8'h33;
			13'h09a0: data_buf = 8'hc5;
			13'h09a1: data_buf = 8'hcd;
			13'h09a2: data_buf = 8'h19;
			13'h09a3: data_buf = 8'h09;
			13'h09a4: data_buf = 8'hcd;
			13'h09a5: data_buf = 8'he6;
			13'h09a6: data_buf = 8'h09;
			13'h09a7: data_buf = 8'he5;
			13'h09a8: data_buf = 8'h2a;
			13'h09a9: data_buf = 8'ha1;
			13'h09aa: data_buf = 8'h80;
			13'h09ab: data_buf = 8'hcd;
			13'h09ac: data_buf = 8'hbd;
			13'h09ad: data_buf = 8'h06;
			13'h09ae: data_buf = 8'he1;
			13'h09af: data_buf = 8'h23;
			13'h09b0: data_buf = 8'hdc;
			13'h09b1: data_buf = 8'he4;
			13'h09b2: data_buf = 8'h04;
			13'h09b3: data_buf = 8'hd4;
			13'h09b4: data_buf = 8'he1;
			13'h09b5: data_buf = 8'h04;
			13'h09b6: data_buf = 8'h60;
			13'h09b7: data_buf = 8'h69;
			13'h09b8: data_buf = 8'h2b;
			13'h09b9: data_buf = 8'hd8;
			13'h09ba: data_buf = 8'h1e;
			13'h09bb: data_buf = 8'h0e;
			13'h09bc: data_buf = 8'hc3;
			13'h09bd: data_buf = 8'h09;
			13'h09be: data_buf = 8'h04;
			13'h09bf: data_buf = 8'hc0;
			13'h09c0: data_buf = 8'h16;
			13'h09c1: data_buf = 8'hff;
			13'h09c2: data_buf = 8'hcd;
			13'h09c3: data_buf = 8'h9e;
			13'h09c4: data_buf = 8'h03;
			13'h09c5: data_buf = 8'hf9;
			13'h09c6: data_buf = 8'hfe;
			13'h09c7: data_buf = 8'h8c;
			13'h09c8: data_buf = 8'h1e;
			13'h09c9: data_buf = 8'h04;
			13'h09ca: data_buf = 8'hc2;
			13'h09cb: data_buf = 8'h09;
			13'h09cc: data_buf = 8'h04;
			13'h09cd: data_buf = 8'he1;
			13'h09ce: data_buf = 8'h22;
			13'h09cf: data_buf = 8'ha1;
			13'h09d0: data_buf = 8'h80;
			13'h09d1: data_buf = 8'h23;
			13'h09d2: data_buf = 8'h7c;
			13'h09d3: data_buf = 8'hb5;
			13'h09d4: data_buf = 8'hc2;
			13'h09d5: data_buf = 8'hde;
			13'h09d6: data_buf = 8'h09;
			13'h09d7: data_buf = 8'h3a;
			13'h09d8: data_buf = 8'h11;
			13'h09d9: data_buf = 8'h81;
			13'h09da: data_buf = 8'hb7;
			13'h09db: data_buf = 8'hc2;
			13'h09dc: data_buf = 8'h3f;
			13'h09dd: data_buf = 8'h04;
			13'h09de: data_buf = 8'h21;
			13'h09df: data_buf = 8'h0d;
			13'h09e0: data_buf = 8'h08;
			13'h09e1: data_buf = 8'he3;
			13'h09e2: data_buf = 8'h3e;
			13'h09e3: data_buf = 8'he1;
			13'h09e4: data_buf = 8'h01;
			13'h09e5: data_buf = 8'h3a;
			13'h09e6: data_buf = 8'h0e;
			13'h09e7: data_buf = 8'h00;
			13'h09e8: data_buf = 8'h06;
			13'h09e9: data_buf = 8'h00;
			13'h09ea: data_buf = 8'h79;
			13'h09eb: data_buf = 8'h48;
			13'h09ec: data_buf = 8'h47;
			13'h09ed: data_buf = 8'h7e;
			13'h09ee: data_buf = 8'hb7;
			13'h09ef: data_buf = 8'hc8;
			13'h09f0: data_buf = 8'hb8;
			13'h09f1: data_buf = 8'hc8;
			13'h09f2: data_buf = 8'h23;
			13'h09f3: data_buf = 8'hfe;
			13'h09f4: data_buf = 8'h22;
			13'h09f5: data_buf = 8'hca;
			13'h09f6: data_buf = 8'hea;
			13'h09f7: data_buf = 8'h09;
			13'h09f8: data_buf = 8'hc3;
			13'h09f9: data_buf = 8'hed;
			13'h09fa: data_buf = 8'h09;
			13'h09fb: data_buf = 8'hcd;
			13'h09fc: data_buf = 8'hb0;
			13'h09fd: data_buf = 8'h0e;
			13'h09fe: data_buf = 8'hcd;
			13'h09ff: data_buf = 8'hc3;
			13'h0a00: data_buf = 8'h06;
			13'h0a01: data_buf = 8'hb4;
			13'h0a02: data_buf = 8'hd5;
			13'h0a03: data_buf = 8'h3a;
			13'h0a04: data_buf = 8'hf2;
			13'h0a05: data_buf = 8'h80;
			13'h0a06: data_buf = 8'hf5;
			13'h0a07: data_buf = 8'hcd;
			13'h0a08: data_buf = 8'hcc;
			13'h0a09: data_buf = 8'h0c;
			13'h0a0a: data_buf = 8'hf1;
			13'h0a0b: data_buf = 8'he3;
			13'h0a0c: data_buf = 8'h22;
			13'h0a0d: data_buf = 8'h13;
			13'h0a0e: data_buf = 8'h81;
			13'h0a0f: data_buf = 8'h1f;
			13'h0a10: data_buf = 8'hcd;
			13'h0a11: data_buf = 8'hbf;
			13'h0a12: data_buf = 8'h0c;
			13'h0a13: data_buf = 8'hca;
			13'h0a14: data_buf = 8'h4e;
			13'h0a15: data_buf = 8'h0a;
			13'h0a16: data_buf = 8'he5;
			13'h0a17: data_buf = 8'h2a;
			13'h0a18: data_buf = 8'h29;
			13'h0a19: data_buf = 8'h81;
			13'h0a1a: data_buf = 8'he5;
			13'h0a1b: data_buf = 8'h23;
			13'h0a1c: data_buf = 8'h23;
			13'h0a1d: data_buf = 8'h5e;
			13'h0a1e: data_buf = 8'h23;
			13'h0a1f: data_buf = 8'h56;
			13'h0a20: data_buf = 8'h2a;
			13'h0a21: data_buf = 8'ha3;
			13'h0a22: data_buf = 8'h80;
			13'h0a23: data_buf = 8'hcd;
			13'h0a24: data_buf = 8'hbd;
			13'h0a25: data_buf = 8'h06;
			13'h0a26: data_buf = 8'hd2;
			13'h0a27: data_buf = 8'h3d;
			13'h0a28: data_buf = 8'h0a;
			13'h0a29: data_buf = 8'h2a;
			13'h0a2a: data_buf = 8'h9f;
			13'h0a2b: data_buf = 8'h80;
			13'h0a2c: data_buf = 8'hcd;
			13'h0a2d: data_buf = 8'hbd;
			13'h0a2e: data_buf = 8'h06;
			13'h0a2f: data_buf = 8'hd1;
			13'h0a30: data_buf = 8'hd2;
			13'h0a31: data_buf = 8'h45;
			13'h0a32: data_buf = 8'h0a;
			13'h0a33: data_buf = 8'h21;
			13'h0a34: data_buf = 8'h04;
			13'h0a35: data_buf = 8'h81;
			13'h0a36: data_buf = 8'hcd;
			13'h0a37: data_buf = 8'hbd;
			13'h0a38: data_buf = 8'h06;
			13'h0a39: data_buf = 8'hd2;
			13'h0a3a: data_buf = 8'h45;
			13'h0a3b: data_buf = 8'h0a;
			13'h0a3c: data_buf = 8'h3e;
			13'h0a3d: data_buf = 8'hd1;
			13'h0a3e: data_buf = 8'hcd;
			13'h0a3f: data_buf = 8'hf4;
			13'h0a40: data_buf = 8'h12;
			13'h0a41: data_buf = 8'heb;
			13'h0a42: data_buf = 8'hcd;
			13'h0a43: data_buf = 8'h2d;
			13'h0a44: data_buf = 8'h11;
			13'h0a45: data_buf = 8'hcd;
			13'h0a46: data_buf = 8'hf4;
			13'h0a47: data_buf = 8'h12;
			13'h0a48: data_buf = 8'he1;
			13'h0a49: data_buf = 8'hcd;
			13'h0a4a: data_buf = 8'hf7;
			13'h0a4b: data_buf = 8'h16;
			13'h0a4c: data_buf = 8'he1;
			13'h0a4d: data_buf = 8'hc9;
			13'h0a4e: data_buf = 8'he5;
			13'h0a4f: data_buf = 8'hcd;
			13'h0a50: data_buf = 8'hf4;
			13'h0a51: data_buf = 8'h16;
			13'h0a52: data_buf = 8'hd1;
			13'h0a53: data_buf = 8'he1;
			13'h0a54: data_buf = 8'hc9;
			13'h0a55: data_buf = 8'hcd;
			13'h0a56: data_buf = 8'h1b;
			13'h0a57: data_buf = 8'h14;
			13'h0a58: data_buf = 8'h7e;
			13'h0a59: data_buf = 8'h47;
			13'h0a5a: data_buf = 8'hfe;
			13'h0a5b: data_buf = 8'h8c;
			13'h0a5c: data_buf = 8'hca;
			13'h0a5d: data_buf = 8'h64;
			13'h0a5e: data_buf = 8'h0a;
			13'h0a5f: data_buf = 8'hcd;
			13'h0a60: data_buf = 8'hc3;
			13'h0a61: data_buf = 8'h06;
			13'h0a62: data_buf = 8'h88;
			13'h0a63: data_buf = 8'h2b;
			13'h0a64: data_buf = 8'h4b;
			13'h0a65: data_buf = 8'h0d;
			13'h0a66: data_buf = 8'h78;
			13'h0a67: data_buf = 8'hca;
			13'h0a68: data_buf = 8'h35;
			13'h0a69: data_buf = 8'h08;
			13'h0a6a: data_buf = 8'hcd;
			13'h0a6b: data_buf = 8'h1a;
			13'h0a6c: data_buf = 8'h09;
			13'h0a6d: data_buf = 8'hfe;
			13'h0a6e: data_buf = 8'h2c;
			13'h0a6f: data_buf = 8'hc0;
			13'h0a70: data_buf = 8'hc3;
			13'h0a71: data_buf = 8'h65;
			13'h0a72: data_buf = 8'h0a;
			13'h0a73: data_buf = 8'hcd;
			13'h0a74: data_buf = 8'hcc;
			13'h0a75: data_buf = 8'h0c;
			13'h0a76: data_buf = 8'h7e;
			13'h0a77: data_buf = 8'hfe;
			13'h0a78: data_buf = 8'h88;
			13'h0a79: data_buf = 8'hca;
			13'h0a7a: data_buf = 8'h81;
			13'h0a7b: data_buf = 8'h0a;
			13'h0a7c: data_buf = 8'hcd;
			13'h0a7d: data_buf = 8'hc3;
			13'h0a7e: data_buf = 8'h06;
			13'h0a7f: data_buf = 8'ha9;
			13'h0a80: data_buf = 8'h2b;
			13'h0a81: data_buf = 8'hcd;
			13'h0a82: data_buf = 8'hbd;
			13'h0a83: data_buf = 8'h0c;
			13'h0a84: data_buf = 8'hcd;
			13'h0a85: data_buf = 8'h9c;
			13'h0a86: data_buf = 8'h16;
			13'h0a87: data_buf = 8'hca;
			13'h0a88: data_buf = 8'he6;
			13'h0a89: data_buf = 8'h09;
			13'h0a8a: data_buf = 8'hcd;
			13'h0a8b: data_buf = 8'h4d;
			13'h0a8c: data_buf = 8'h08;
			13'h0a8d: data_buf = 8'hda;
			13'h0a8e: data_buf = 8'ha1;
			13'h0a8f: data_buf = 8'h09;
			13'h0a90: data_buf = 8'hc3;
			13'h0a91: data_buf = 8'h34;
			13'h0a92: data_buf = 8'h08;
			13'h0a93: data_buf = 8'h2b;
			13'h0a94: data_buf = 8'hcd;
			13'h0a95: data_buf = 8'h4d;
			13'h0a96: data_buf = 8'h08;
			13'h0a97: data_buf = 8'hca;
			13'h0a98: data_buf = 8'hf5;
			13'h0a99: data_buf = 8'h0a;
			13'h0a9a: data_buf = 8'hc8;
			13'h0a9b: data_buf = 8'hfe;
			13'h0a9c: data_buf = 8'ha5;
			13'h0a9d: data_buf = 8'hca;
			13'h0a9e: data_buf = 8'h28;
			13'h0a9f: data_buf = 8'h0b;
			13'h0aa0: data_buf = 8'hfe;
			13'h0aa1: data_buf = 8'ha8;
			13'h0aa2: data_buf = 8'hca;
			13'h0aa3: data_buf = 8'h28;
			13'h0aa4: data_buf = 8'h0b;
			13'h0aa5: data_buf = 8'he5;
			13'h0aa6: data_buf = 8'hfe;
			13'h0aa7: data_buf = 8'h2c;
			13'h0aa8: data_buf = 8'hca;
			13'h0aa9: data_buf = 8'h11;
			13'h0aaa: data_buf = 8'h0b;
			13'h0aab: data_buf = 8'hfe;
			13'h0aac: data_buf = 8'h3b;
			13'h0aad: data_buf = 8'hca;
			13'h0aae: data_buf = 8'h4b;
			13'h0aaf: data_buf = 8'h0b;
			13'h0ab0: data_buf = 8'hc1;
			13'h0ab1: data_buf = 8'hcd;
			13'h0ab2: data_buf = 8'hcc;
			13'h0ab3: data_buf = 8'h0c;
			13'h0ab4: data_buf = 8'he5;
			13'h0ab5: data_buf = 8'h3a;
			13'h0ab6: data_buf = 8'hf2;
			13'h0ab7: data_buf = 8'h80;
			13'h0ab8: data_buf = 8'hb7;
			13'h0ab9: data_buf = 8'hc2;
			13'h0aba: data_buf = 8'he1;
			13'h0abb: data_buf = 8'h0a;
			13'h0abc: data_buf = 8'hcd;
			13'h0abd: data_buf = 8'h41;
			13'h0abe: data_buf = 8'h18;
			13'h0abf: data_buf = 8'hcd;
			13'h0ac0: data_buf = 8'h51;
			13'h0ac1: data_buf = 8'h11;
			13'h0ac2: data_buf = 8'h36;
			13'h0ac3: data_buf = 8'h20;
			13'h0ac4: data_buf = 8'h2a;
			13'h0ac5: data_buf = 8'h29;
			13'h0ac6: data_buf = 8'h81;
			13'h0ac7: data_buf = 8'h34;
			13'h0ac8: data_buf = 8'h2a;
			13'h0ac9: data_buf = 8'h29;
			13'h0aca: data_buf = 8'h81;
			13'h0acb: data_buf = 8'h3a;
			13'h0acc: data_buf = 8'h87;
			13'h0acd: data_buf = 8'h80;
			13'h0ace: data_buf = 8'h47;
			13'h0acf: data_buf = 8'h04;
			13'h0ad0: data_buf = 8'hca;
			13'h0ad1: data_buf = 8'hdd;
			13'h0ad2: data_buf = 8'h0a;
			13'h0ad3: data_buf = 8'h04;
			13'h0ad4: data_buf = 8'h3a;
			13'h0ad5: data_buf = 8'hf0;
			13'h0ad6: data_buf = 8'h80;
			13'h0ad7: data_buf = 8'h86;
			13'h0ad8: data_buf = 8'h3d;
			13'h0ad9: data_buf = 8'hb8;
			13'h0ada: data_buf = 8'hd4;
			13'h0adb: data_buf = 8'hf5;
			13'h0adc: data_buf = 8'h0a;
			13'h0add: data_buf = 8'hcd;
			13'h0ade: data_buf = 8'h96;
			13'h0adf: data_buf = 8'h11;
			13'h0ae0: data_buf = 8'haf;
			13'h0ae1: data_buf = 8'hc4;
			13'h0ae2: data_buf = 8'h96;
			13'h0ae3: data_buf = 8'h11;
			13'h0ae4: data_buf = 8'he1;
			13'h0ae5: data_buf = 8'hc3;
			13'h0ae6: data_buf = 8'h93;
			13'h0ae7: data_buf = 8'h0a;
			13'h0ae8: data_buf = 8'h3a;
			13'h0ae9: data_buf = 8'hf0;
			13'h0aea: data_buf = 8'h80;
			13'h0aeb: data_buf = 8'hb7;
			13'h0aec: data_buf = 8'hc8;
			13'h0aed: data_buf = 8'hc3;
			13'h0aee: data_buf = 8'hf5;
			13'h0aef: data_buf = 8'h0a;
			13'h0af0: data_buf = 8'h36;
			13'h0af1: data_buf = 8'h00;
			13'h0af2: data_buf = 8'h21;
			13'h0af3: data_buf = 8'ha5;
			13'h0af4: data_buf = 8'h80;
			13'h0af5: data_buf = 8'h3e;
			13'h0af6: data_buf = 8'h0d;
			13'h0af7: data_buf = 8'hcd;
			13'h0af8: data_buf = 8'hce;
			13'h0af9: data_buf = 8'h06;
			13'h0afa: data_buf = 8'h3e;
			13'h0afb: data_buf = 8'h0a;
			13'h0afc: data_buf = 8'hcd;
			13'h0afd: data_buf = 8'hce;
			13'h0afe: data_buf = 8'h06;
			13'h0aff: data_buf = 8'haf;
			13'h0b00: data_buf = 8'h32;
			13'h0b01: data_buf = 8'hf0;
			13'h0b02: data_buf = 8'h80;
			13'h0b03: data_buf = 8'h3a;
			13'h0b04: data_buf = 8'h86;
			13'h0b05: data_buf = 8'h80;
			13'h0b06: data_buf = 8'h3d;
			13'h0b07: data_buf = 8'hc8;
			13'h0b08: data_buf = 8'hf5;
			13'h0b09: data_buf = 8'haf;
			13'h0b0a: data_buf = 8'hcd;
			13'h0b0b: data_buf = 8'hce;
			13'h0b0c: data_buf = 8'h06;
			13'h0b0d: data_buf = 8'hf1;
			13'h0b0e: data_buf = 8'hc3;
			13'h0b0f: data_buf = 8'h06;
			13'h0b10: data_buf = 8'h0b;
			13'h0b11: data_buf = 8'h3a;
			13'h0b12: data_buf = 8'h88;
			13'h0b13: data_buf = 8'h80;
			13'h0b14: data_buf = 8'h47;
			13'h0b15: data_buf = 8'h3a;
			13'h0b16: data_buf = 8'hf0;
			13'h0b17: data_buf = 8'h80;
			13'h0b18: data_buf = 8'hb8;
			13'h0b19: data_buf = 8'hd4;
			13'h0b1a: data_buf = 8'hf5;
			13'h0b1b: data_buf = 8'h0a;
			13'h0b1c: data_buf = 8'hd2;
			13'h0b1d: data_buf = 8'h4b;
			13'h0b1e: data_buf = 8'h0b;
			13'h0b1f: data_buf = 8'hd6;
			13'h0b20: data_buf = 8'h0e;
			13'h0b21: data_buf = 8'hd2;
			13'h0b22: data_buf = 8'h1f;
			13'h0b23: data_buf = 8'h0b;
			13'h0b24: data_buf = 8'h2f;
			13'h0b25: data_buf = 8'hc3;
			13'h0b26: data_buf = 8'h40;
			13'h0b27: data_buf = 8'h0b;
			13'h0b28: data_buf = 8'hf5;
			13'h0b29: data_buf = 8'hcd;
			13'h0b2a: data_buf = 8'h18;
			13'h0b2b: data_buf = 8'h14;
			13'h0b2c: data_buf = 8'hcd;
			13'h0b2d: data_buf = 8'hc3;
			13'h0b2e: data_buf = 8'h06;
			13'h0b2f: data_buf = 8'h29;
			13'h0b30: data_buf = 8'h2b;
			13'h0b31: data_buf = 8'hf1;
			13'h0b32: data_buf = 8'hd6;
			13'h0b33: data_buf = 8'ha8;
			13'h0b34: data_buf = 8'he5;
			13'h0b35: data_buf = 8'hca;
			13'h0b36: data_buf = 8'h3b;
			13'h0b37: data_buf = 8'h0b;
			13'h0b38: data_buf = 8'h3a;
			13'h0b39: data_buf = 8'hf0;
			13'h0b3a: data_buf = 8'h80;
			13'h0b3b: data_buf = 8'h2f;
			13'h0b3c: data_buf = 8'h83;
			13'h0b3d: data_buf = 8'hd2;
			13'h0b3e: data_buf = 8'h4b;
			13'h0b3f: data_buf = 8'h0b;
			13'h0b40: data_buf = 8'h3c;
			13'h0b41: data_buf = 8'h47;
			13'h0b42: data_buf = 8'h3e;
			13'h0b43: data_buf = 8'h20;
			13'h0b44: data_buf = 8'hcd;
			13'h0b45: data_buf = 8'hce;
			13'h0b46: data_buf = 8'h06;
			13'h0b47: data_buf = 8'h05;
			13'h0b48: data_buf = 8'hc2;
			13'h0b49: data_buf = 8'h44;
			13'h0b4a: data_buf = 8'h0b;
			13'h0b4b: data_buf = 8'he1;
			13'h0b4c: data_buf = 8'hcd;
			13'h0b4d: data_buf = 8'h4d;
			13'h0b4e: data_buf = 8'h08;
			13'h0b4f: data_buf = 8'hc3;
			13'h0b50: data_buf = 8'h9a;
			13'h0b51: data_buf = 8'h0a;
			13'h0b52: data_buf = 8'h3f;
			13'h0b53: data_buf = 8'h52;
			13'h0b54: data_buf = 8'h65;
			13'h0b55: data_buf = 8'h64;
			13'h0b56: data_buf = 8'h6f;
			13'h0b57: data_buf = 8'h20;
			13'h0b58: data_buf = 8'h66;
			13'h0b59: data_buf = 8'h72;
			13'h0b5a: data_buf = 8'h6f;
			13'h0b5b: data_buf = 8'h6d;
			13'h0b5c: data_buf = 8'h20;
			13'h0b5d: data_buf = 8'h73;
			13'h0b5e: data_buf = 8'h74;
			13'h0b5f: data_buf = 8'h61;
			13'h0b60: data_buf = 8'h72;
			13'h0b61: data_buf = 8'h74;
			13'h0b62: data_buf = 8'h0d;
			13'h0b63: data_buf = 8'h0a;
			13'h0b64: data_buf = 8'h00;
			13'h0b65: data_buf = 8'h3a;
			13'h0b66: data_buf = 8'h12;
			13'h0b67: data_buf = 8'h81;
			13'h0b68: data_buf = 8'hb7;
			13'h0b69: data_buf = 8'hc2;
			13'h0b6a: data_buf = 8'hef;
			13'h0b6b: data_buf = 8'h03;
			13'h0b6c: data_buf = 8'hc1;
			13'h0b6d: data_buf = 8'h21;
			13'h0b6e: data_buf = 8'h52;
			13'h0b6f: data_buf = 8'h0b;
			13'h0b70: data_buf = 8'hcd;
			13'h0b71: data_buf = 8'h93;
			13'h0b72: data_buf = 8'h11;
			13'h0b73: data_buf = 8'hc3;
			13'h0b74: data_buf = 8'h40;
			13'h0b75: data_buf = 8'h05;
			13'h0b76: data_buf = 8'hcd;
			13'h0b77: data_buf = 8'hfe;
			13'h0b78: data_buf = 8'h10;
			13'h0b79: data_buf = 8'h7e;
			13'h0b7a: data_buf = 8'hfe;
			13'h0b7b: data_buf = 8'h22;
			13'h0b7c: data_buf = 8'h3e;
			13'h0b7d: data_buf = 8'h00;
			13'h0b7e: data_buf = 8'h32;
			13'h0b7f: data_buf = 8'h8a;
			13'h0b80: data_buf = 8'h80;
			13'h0b81: data_buf = 8'hc2;
			13'h0b82: data_buf = 8'h90;
			13'h0b83: data_buf = 8'h0b;
			13'h0b84: data_buf = 8'hcd;
			13'h0b85: data_buf = 8'h52;
			13'h0b86: data_buf = 8'h11;
			13'h0b87: data_buf = 8'hcd;
			13'h0b88: data_buf = 8'hc3;
			13'h0b89: data_buf = 8'h06;
			13'h0b8a: data_buf = 8'h3b;
			13'h0b8b: data_buf = 8'he5;
			13'h0b8c: data_buf = 8'hcd;
			13'h0b8d: data_buf = 8'h96;
			13'h0b8e: data_buf = 8'h11;
			13'h0b8f: data_buf = 8'h3e;
			13'h0b90: data_buf = 8'he5;
			13'h0b91: data_buf = 8'hcd;
			13'h0b92: data_buf = 8'h44;
			13'h0b93: data_buf = 8'h05;
			13'h0b94: data_buf = 8'hc1;
			13'h0b95: data_buf = 8'hda;
			13'h0b96: data_buf = 8'h9c;
			13'h0b97: data_buf = 8'h08;
			13'h0b98: data_buf = 8'h23;
			13'h0b99: data_buf = 8'h7e;
			13'h0b9a: data_buf = 8'hb7;
			13'h0b9b: data_buf = 8'h2b;
			13'h0b9c: data_buf = 8'hc5;
			13'h0b9d: data_buf = 8'hca;
			13'h0b9e: data_buf = 8'he3;
			13'h0b9f: data_buf = 8'h09;
			13'h0ba0: data_buf = 8'h36;
			13'h0ba1: data_buf = 8'h2c;
			13'h0ba2: data_buf = 8'hc3;
			13'h0ba3: data_buf = 8'haa;
			13'h0ba4: data_buf = 8'h0b;
			13'h0ba5: data_buf = 8'he5;
			13'h0ba6: data_buf = 8'h2a;
			13'h0ba7: data_buf = 8'h21;
			13'h0ba8: data_buf = 8'h81;
			13'h0ba9: data_buf = 8'hf6;
			13'h0baa: data_buf = 8'haf;
			13'h0bab: data_buf = 8'h32;
			13'h0bac: data_buf = 8'h12;
			13'h0bad: data_buf = 8'h81;
			13'h0bae: data_buf = 8'he3;
			13'h0baf: data_buf = 8'hc3;
			13'h0bb0: data_buf = 8'hb6;
			13'h0bb1: data_buf = 8'h0b;
			13'h0bb2: data_buf = 8'hcd;
			13'h0bb3: data_buf = 8'hc3;
			13'h0bb4: data_buf = 8'h06;
			13'h0bb5: data_buf = 8'h2c;
			13'h0bb6: data_buf = 8'hcd;
			13'h0bb7: data_buf = 8'hb0;
			13'h0bb8: data_buf = 8'h0e;
			13'h0bb9: data_buf = 8'he3;
			13'h0bba: data_buf = 8'hd5;
			13'h0bbb: data_buf = 8'h7e;
			13'h0bbc: data_buf = 8'hfe;
			13'h0bbd: data_buf = 8'h2c;
			13'h0bbe: data_buf = 8'hca;
			13'h0bbf: data_buf = 8'hde;
			13'h0bc0: data_buf = 8'h0b;
			13'h0bc1: data_buf = 8'h3a;
			13'h0bc2: data_buf = 8'h12;
			13'h0bc3: data_buf = 8'h81;
			13'h0bc4: data_buf = 8'hb7;
			13'h0bc5: data_buf = 8'hc2;
			13'h0bc6: data_buf = 8'h4b;
			13'h0bc7: data_buf = 8'h0c;
			13'h0bc8: data_buf = 8'h3e;
			13'h0bc9: data_buf = 8'h3f;
			13'h0bca: data_buf = 8'hcd;
			13'h0bcb: data_buf = 8'hce;
			13'h0bcc: data_buf = 8'h06;
			13'h0bcd: data_buf = 8'hcd;
			13'h0bce: data_buf = 8'h44;
			13'h0bcf: data_buf = 8'h05;
			13'h0bd0: data_buf = 8'hd1;
			13'h0bd1: data_buf = 8'hc1;
			13'h0bd2: data_buf = 8'hda;
			13'h0bd3: data_buf = 8'h9c;
			13'h0bd4: data_buf = 8'h08;
			13'h0bd5: data_buf = 8'h23;
			13'h0bd6: data_buf = 8'h7e;
			13'h0bd7: data_buf = 8'hb7;
			13'h0bd8: data_buf = 8'h2b;
			13'h0bd9: data_buf = 8'hc5;
			13'h0bda: data_buf = 8'hca;
			13'h0bdb: data_buf = 8'he3;
			13'h0bdc: data_buf = 8'h09;
			13'h0bdd: data_buf = 8'hd5;
			13'h0bde: data_buf = 8'h3a;
			13'h0bdf: data_buf = 8'hf2;
			13'h0be0: data_buf = 8'h80;
			13'h0be1: data_buf = 8'hb7;
			13'h0be2: data_buf = 8'hca;
			13'h0be3: data_buf = 8'h08;
			13'h0be4: data_buf = 8'h0c;
			13'h0be5: data_buf = 8'hcd;
			13'h0be6: data_buf = 8'h4d;
			13'h0be7: data_buf = 8'h08;
			13'h0be8: data_buf = 8'h57;
			13'h0be9: data_buf = 8'h47;
			13'h0bea: data_buf = 8'hfe;
			13'h0beb: data_buf = 8'h22;
			13'h0bec: data_buf = 8'hca;
			13'h0bed: data_buf = 8'hfc;
			13'h0bee: data_buf = 8'h0b;
			13'h0bef: data_buf = 8'h3a;
			13'h0bf0: data_buf = 8'h12;
			13'h0bf1: data_buf = 8'h81;
			13'h0bf2: data_buf = 8'hb7;
			13'h0bf3: data_buf = 8'h57;
			13'h0bf4: data_buf = 8'hca;
			13'h0bf5: data_buf = 8'hf9;
			13'h0bf6: data_buf = 8'h0b;
			13'h0bf7: data_buf = 8'h16;
			13'h0bf8: data_buf = 8'h3a;
			13'h0bf9: data_buf = 8'h06;
			13'h0bfa: data_buf = 8'h2c;
			13'h0bfb: data_buf = 8'h2b;
			13'h0bfc: data_buf = 8'hcd;
			13'h0bfd: data_buf = 8'h55;
			13'h0bfe: data_buf = 8'h11;
			13'h0bff: data_buf = 8'heb;
			13'h0c00: data_buf = 8'h21;
			13'h0c01: data_buf = 8'h13;
			13'h0c02: data_buf = 8'h0c;
			13'h0c03: data_buf = 8'he3;
			13'h0c04: data_buf = 8'hd5;
			13'h0c05: data_buf = 8'hc3;
			13'h0c06: data_buf = 8'h16;
			13'h0c07: data_buf = 8'h0a;
			13'h0c08: data_buf = 8'hcd;
			13'h0c09: data_buf = 8'h4d;
			13'h0c0a: data_buf = 8'h08;
			13'h0c0b: data_buf = 8'hcd;
			13'h0c0c: data_buf = 8'ha3;
			13'h0c0d: data_buf = 8'h17;
			13'h0c0e: data_buf = 8'he3;
			13'h0c0f: data_buf = 8'hcd;
			13'h0c10: data_buf = 8'hf4;
			13'h0c11: data_buf = 8'h16;
			13'h0c12: data_buf = 8'he1;
			13'h0c13: data_buf = 8'h2b;
			13'h0c14: data_buf = 8'hcd;
			13'h0c15: data_buf = 8'h4d;
			13'h0c16: data_buf = 8'h08;
			13'h0c17: data_buf = 8'hca;
			13'h0c18: data_buf = 8'h1f;
			13'h0c19: data_buf = 8'h0c;
			13'h0c1a: data_buf = 8'hfe;
			13'h0c1b: data_buf = 8'h2c;
			13'h0c1c: data_buf = 8'hc2;
			13'h0c1d: data_buf = 8'h65;
			13'h0c1e: data_buf = 8'h0b;
			13'h0c1f: data_buf = 8'he3;
			13'h0c20: data_buf = 8'h2b;
			13'h0c21: data_buf = 8'hcd;
			13'h0c22: data_buf = 8'h4d;
			13'h0c23: data_buf = 8'h08;
			13'h0c24: data_buf = 8'hc2;
			13'h0c25: data_buf = 8'hb2;
			13'h0c26: data_buf = 8'h0b;
			13'h0c27: data_buf = 8'hd1;
			13'h0c28: data_buf = 8'h3a;
			13'h0c29: data_buf = 8'h12;
			13'h0c2a: data_buf = 8'h81;
			13'h0c2b: data_buf = 8'hb7;
			13'h0c2c: data_buf = 8'heb;
			13'h0c2d: data_buf = 8'hc2;
			13'h0c2e: data_buf = 8'h73;
			13'h0c2f: data_buf = 8'h08;
			13'h0c30: data_buf = 8'hd5;
			13'h0c31: data_buf = 8'hb6;
			13'h0c32: data_buf = 8'h21;
			13'h0c33: data_buf = 8'h3a;
			13'h0c34: data_buf = 8'h0c;
			13'h0c35: data_buf = 8'hc4;
			13'h0c36: data_buf = 8'h93;
			13'h0c37: data_buf = 8'h11;
			13'h0c38: data_buf = 8'he1;
			13'h0c39: data_buf = 8'hc9;
			13'h0c3a: data_buf = 8'h3f;
			13'h0c3b: data_buf = 8'h45;
			13'h0c3c: data_buf = 8'h78;
			13'h0c3d: data_buf = 8'h74;
			13'h0c3e: data_buf = 8'h72;
			13'h0c3f: data_buf = 8'h61;
			13'h0c40: data_buf = 8'h20;
			13'h0c41: data_buf = 8'h69;
			13'h0c42: data_buf = 8'h67;
			13'h0c43: data_buf = 8'h6e;
			13'h0c44: data_buf = 8'h6f;
			13'h0c45: data_buf = 8'h72;
			13'h0c46: data_buf = 8'h65;
			13'h0c47: data_buf = 8'h64;
			13'h0c48: data_buf = 8'h0d;
			13'h0c49: data_buf = 8'h0a;
			13'h0c4a: data_buf = 8'h00;
			13'h0c4b: data_buf = 8'hcd;
			13'h0c4c: data_buf = 8'he4;
			13'h0c4d: data_buf = 8'h09;
			13'h0c4e: data_buf = 8'hb7;
			13'h0c4f: data_buf = 8'hc2;
			13'h0c50: data_buf = 8'h64;
			13'h0c51: data_buf = 8'h0c;
			13'h0c52: data_buf = 8'h23;
			13'h0c53: data_buf = 8'h7e;
			13'h0c54: data_buf = 8'h23;
			13'h0c55: data_buf = 8'hb6;
			13'h0c56: data_buf = 8'h1e;
			13'h0c57: data_buf = 8'h06;
			13'h0c58: data_buf = 8'hca;
			13'h0c59: data_buf = 8'h09;
			13'h0c5a: data_buf = 8'h04;
			13'h0c5b: data_buf = 8'h23;
			13'h0c5c: data_buf = 8'h5e;
			13'h0c5d: data_buf = 8'h23;
			13'h0c5e: data_buf = 8'h56;
			13'h0c5f: data_buf = 8'heb;
			13'h0c60: data_buf = 8'h22;
			13'h0c61: data_buf = 8'h0e;
			13'h0c62: data_buf = 8'h81;
			13'h0c63: data_buf = 8'heb;
			13'h0c64: data_buf = 8'hcd;
			13'h0c65: data_buf = 8'h4d;
			13'h0c66: data_buf = 8'h08;
			13'h0c67: data_buf = 8'hfe;
			13'h0c68: data_buf = 8'h83;
			13'h0c69: data_buf = 8'hc2;
			13'h0c6a: data_buf = 8'h4b;
			13'h0c6b: data_buf = 8'h0c;
			13'h0c6c: data_buf = 8'hc3;
			13'h0c6d: data_buf = 8'hde;
			13'h0c6e: data_buf = 8'h0b;
			13'h0c6f: data_buf = 8'h11;
			13'h0c70: data_buf = 8'h00;
			13'h0c71: data_buf = 8'h00;
			13'h0c72: data_buf = 8'hc4;
			13'h0c73: data_buf = 8'hb0;
			13'h0c74: data_buf = 8'h0e;
			13'h0c75: data_buf = 8'h22;
			13'h0c76: data_buf = 8'h13;
			13'h0c77: data_buf = 8'h81;
			13'h0c78: data_buf = 8'hcd;
			13'h0c79: data_buf = 8'h9e;
			13'h0c7a: data_buf = 8'h03;
			13'h0c7b: data_buf = 8'hc2;
			13'h0c7c: data_buf = 8'hfb;
			13'h0c7d: data_buf = 8'h03;
			13'h0c7e: data_buf = 8'hf9;
			13'h0c7f: data_buf = 8'hd5;
			13'h0c80: data_buf = 8'h7e;
			13'h0c81: data_buf = 8'h23;
			13'h0c82: data_buf = 8'hf5;
			13'h0c83: data_buf = 8'hd5;
			13'h0c84: data_buf = 8'hcd;
			13'h0c85: data_buf = 8'hda;
			13'h0c86: data_buf = 8'h16;
			13'h0c87: data_buf = 8'he3;
			13'h0c88: data_buf = 8'he5;
			13'h0c89: data_buf = 8'hcd;
			13'h0c8a: data_buf = 8'h47;
			13'h0c8b: data_buf = 8'h14;
			13'h0c8c: data_buf = 8'he1;
			13'h0c8d: data_buf = 8'hcd;
			13'h0c8e: data_buf = 8'hf4;
			13'h0c8f: data_buf = 8'h16;
			13'h0c90: data_buf = 8'he1;
			13'h0c91: data_buf = 8'hcd;
			13'h0c92: data_buf = 8'heb;
			13'h0c93: data_buf = 8'h16;
			13'h0c94: data_buf = 8'he5;
			13'h0c95: data_buf = 8'hcd;
			13'h0c96: data_buf = 8'h17;
			13'h0c97: data_buf = 8'h17;
			13'h0c98: data_buf = 8'he1;
			13'h0c99: data_buf = 8'hc1;
			13'h0c9a: data_buf = 8'h90;
			13'h0c9b: data_buf = 8'hcd;
			13'h0c9c: data_buf = 8'heb;
			13'h0c9d: data_buf = 8'h16;
			13'h0c9e: data_buf = 8'hca;
			13'h0c9f: data_buf = 8'haa;
			13'h0ca0: data_buf = 8'h0c;
			13'h0ca1: data_buf = 8'heb;
			13'h0ca2: data_buf = 8'h22;
			13'h0ca3: data_buf = 8'ha1;
			13'h0ca4: data_buf = 8'h80;
			13'h0ca5: data_buf = 8'h69;
			13'h0ca6: data_buf = 8'h60;
			13'h0ca7: data_buf = 8'hc3;
			13'h0ca8: data_buf = 8'h09;
			13'h0ca9: data_buf = 8'h08;
			13'h0caa: data_buf = 8'hf9;
			13'h0cab: data_buf = 8'h2a;
			13'h0cac: data_buf = 8'h13;
			13'h0cad: data_buf = 8'h81;
			13'h0cae: data_buf = 8'h7e;
			13'h0caf: data_buf = 8'hfe;
			13'h0cb0: data_buf = 8'h2c;
			13'h0cb1: data_buf = 8'hc2;
			13'h0cb2: data_buf = 8'h0d;
			13'h0cb3: data_buf = 8'h08;
			13'h0cb4: data_buf = 8'hcd;
			13'h0cb5: data_buf = 8'h4d;
			13'h0cb6: data_buf = 8'h08;
			13'h0cb7: data_buf = 8'hcd;
			13'h0cb8: data_buf = 8'h72;
			13'h0cb9: data_buf = 8'h0c;
			13'h0cba: data_buf = 8'hcd;
			13'h0cbb: data_buf = 8'hcc;
			13'h0cbc: data_buf = 8'h0c;
			13'h0cbd: data_buf = 8'hf6;
			13'h0cbe: data_buf = 8'h37;
			13'h0cbf: data_buf = 8'h3a;
			13'h0cc0: data_buf = 8'hf2;
			13'h0cc1: data_buf = 8'h80;
			13'h0cc2: data_buf = 8'h8f;
			13'h0cc3: data_buf = 8'hb7;
			13'h0cc4: data_buf = 8'he8;
			13'h0cc5: data_buf = 8'hc3;
			13'h0cc6: data_buf = 8'h07;
			13'h0cc7: data_buf = 8'h04;
			13'h0cc8: data_buf = 8'hcd;
			13'h0cc9: data_buf = 8'hc3;
			13'h0cca: data_buf = 8'h06;
			13'h0ccb: data_buf = 8'h28;
			13'h0ccc: data_buf = 8'h2b;
			13'h0ccd: data_buf = 8'h16;
			13'h0cce: data_buf = 8'h00;
			13'h0ccf: data_buf = 8'hd5;
			13'h0cd0: data_buf = 8'h0e;
			13'h0cd1: data_buf = 8'h01;
			13'h0cd2: data_buf = 8'hcd;
			13'h0cd3: data_buf = 8'hd2;
			13'h0cd4: data_buf = 8'h03;
			13'h0cd5: data_buf = 8'hcd;
			13'h0cd6: data_buf = 8'h43;
			13'h0cd7: data_buf = 8'h0d;
			13'h0cd8: data_buf = 8'h22;
			13'h0cd9: data_buf = 8'h15;
			13'h0cda: data_buf = 8'h81;
			13'h0cdb: data_buf = 8'h2a;
			13'h0cdc: data_buf = 8'h15;
			13'h0cdd: data_buf = 8'h81;
			13'h0cde: data_buf = 8'hc1;
			13'h0cdf: data_buf = 8'h78;
			13'h0ce0: data_buf = 8'hfe;
			13'h0ce1: data_buf = 8'h78;
			13'h0ce2: data_buf = 8'hd4;
			13'h0ce3: data_buf = 8'hbd;
			13'h0ce4: data_buf = 8'h0c;
			13'h0ce5: data_buf = 8'h7e;
			13'h0ce6: data_buf = 8'h16;
			13'h0ce7: data_buf = 8'h00;
			13'h0ce8: data_buf = 8'hd6;
			13'h0ce9: data_buf = 8'hb3;
			13'h0cea: data_buf = 8'hda;
			13'h0ceb: data_buf = 8'h04;
			13'h0cec: data_buf = 8'h0d;
			13'h0ced: data_buf = 8'hfe;
			13'h0cee: data_buf = 8'h03;
			13'h0cef: data_buf = 8'hd2;
			13'h0cf0: data_buf = 8'h04;
			13'h0cf1: data_buf = 8'h0d;
			13'h0cf2: data_buf = 8'hfe;
			13'h0cf3: data_buf = 8'h01;
			13'h0cf4: data_buf = 8'h17;
			13'h0cf5: data_buf = 8'haa;
			13'h0cf6: data_buf = 8'hba;
			13'h0cf7: data_buf = 8'h57;
			13'h0cf8: data_buf = 8'hda;
			13'h0cf9: data_buf = 8'hf5;
			13'h0cfa: data_buf = 8'h03;
			13'h0cfb: data_buf = 8'h22;
			13'h0cfc: data_buf = 8'h0a;
			13'h0cfd: data_buf = 8'h81;
			13'h0cfe: data_buf = 8'hcd;
			13'h0cff: data_buf = 8'h4d;
			13'h0d00: data_buf = 8'h08;
			13'h0d01: data_buf = 8'hc3;
			13'h0d02: data_buf = 8'he8;
			13'h0d03: data_buf = 8'h0c;
			13'h0d04: data_buf = 8'h7a;
			13'h0d05: data_buf = 8'hb7;
			13'h0d06: data_buf = 8'hc2;
			13'h0d07: data_buf = 8'h2b;
			13'h0d08: data_buf = 8'h0e;
			13'h0d09: data_buf = 8'h7e;
			13'h0d0a: data_buf = 8'h22;
			13'h0d0b: data_buf = 8'h0a;
			13'h0d0c: data_buf = 8'h81;
			13'h0d0d: data_buf = 8'hd6;
			13'h0d0e: data_buf = 8'hac;
			13'h0d0f: data_buf = 8'hd8;
			13'h0d10: data_buf = 8'hfe;
			13'h0d11: data_buf = 8'h07;
			13'h0d12: data_buf = 8'hd0;
			13'h0d13: data_buf = 8'h5f;
			13'h0d14: data_buf = 8'h3a;
			13'h0d15: data_buf = 8'hf2;
			13'h0d16: data_buf = 8'h80;
			13'h0d17: data_buf = 8'h3d;
			13'h0d18: data_buf = 8'hb3;
			13'h0d19: data_buf = 8'h7b;
			13'h0d1a: data_buf = 8'hca;
			13'h0d1b: data_buf = 8'h89;
			13'h0d1c: data_buf = 8'h12;
			13'h0d1d: data_buf = 8'h07;
			13'h0d1e: data_buf = 8'h83;
			13'h0d1f: data_buf = 8'h5f;
			13'h0d20: data_buf = 8'h21;
			13'h0d21: data_buf = 8'he7;
			13'h0d22: data_buf = 8'h02;
			13'h0d23: data_buf = 8'h19;
			13'h0d24: data_buf = 8'h78;
			13'h0d25: data_buf = 8'h56;
			13'h0d26: data_buf = 8'hba;
			13'h0d27: data_buf = 8'hd0;
			13'h0d28: data_buf = 8'h23;
			13'h0d29: data_buf = 8'hcd;
			13'h0d2a: data_buf = 8'hbd;
			13'h0d2b: data_buf = 8'h0c;
			13'h0d2c: data_buf = 8'hc5;
			13'h0d2d: data_buf = 8'h01;
			13'h0d2e: data_buf = 8'hdb;
			13'h0d2f: data_buf = 8'h0c;
			13'h0d30: data_buf = 8'hc5;
			13'h0d31: data_buf = 8'h43;
			13'h0d32: data_buf = 8'h4a;
			13'h0d33: data_buf = 8'hcd;
			13'h0d34: data_buf = 8'hcd;
			13'h0d35: data_buf = 8'h16;
			13'h0d36: data_buf = 8'h58;
			13'h0d37: data_buf = 8'h51;
			13'h0d38: data_buf = 8'h4e;
			13'h0d39: data_buf = 8'h23;
			13'h0d3a: data_buf = 8'h46;
			13'h0d3b: data_buf = 8'h23;
			13'h0d3c: data_buf = 8'hc5;
			13'h0d3d: data_buf = 8'h2a;
			13'h0d3e: data_buf = 8'h0a;
			13'h0d3f: data_buf = 8'h81;
			13'h0d40: data_buf = 8'hc3;
			13'h0d41: data_buf = 8'hcf;
			13'h0d42: data_buf = 8'h0c;
			13'h0d43: data_buf = 8'haf;
			13'h0d44: data_buf = 8'h32;
			13'h0d45: data_buf = 8'hf2;
			13'h0d46: data_buf = 8'h80;
			13'h0d47: data_buf = 8'hcd;
			13'h0d48: data_buf = 8'h4d;
			13'h0d49: data_buf = 8'h08;
			13'h0d4a: data_buf = 8'h1e;
			13'h0d4b: data_buf = 8'h24;
			13'h0d4c: data_buf = 8'hca;
			13'h0d4d: data_buf = 8'h09;
			13'h0d4e: data_buf = 8'h04;
			13'h0d4f: data_buf = 8'hda;
			13'h0d50: data_buf = 8'ha3;
			13'h0d51: data_buf = 8'h17;
			13'h0d52: data_buf = 8'hcd;
			13'h0d53: data_buf = 8'heb;
			13'h0d54: data_buf = 8'h08;
			13'h0d55: data_buf = 8'hd2;
			13'h0d56: data_buf = 8'haa;
			13'h0d57: data_buf = 8'h0d;
			13'h0d58: data_buf = 8'hfe;
			13'h0d59: data_buf = 8'h26;
			13'h0d5a: data_buf = 8'h20;
			13'h0d5b: data_buf = 8'h12;
			13'h0d5c: data_buf = 8'hcd;
			13'h0d5d: data_buf = 8'h4d;
			13'h0d5e: data_buf = 8'h08;
			13'h0d5f: data_buf = 8'hfe;
			13'h0d60: data_buf = 8'h48;
			13'h0d61: data_buf = 8'hca;
			13'h0d62: data_buf = 8'he7;
			13'h0d63: data_buf = 8'h1b;
			13'h0d64: data_buf = 8'hfe;
			13'h0d65: data_buf = 8'h42;
			13'h0d66: data_buf = 8'hca;
			13'h0d67: data_buf = 8'h57;
			13'h0d68: data_buf = 8'h1c;
			13'h0d69: data_buf = 8'h1e;
			13'h0d6a: data_buf = 8'h02;
			13'h0d6b: data_buf = 8'hca;
			13'h0d6c: data_buf = 8'h09;
			13'h0d6d: data_buf = 8'h04;
			13'h0d6e: data_buf = 8'hfe;
			13'h0d6f: data_buf = 8'hac;
			13'h0d70: data_buf = 8'hca;
			13'h0d71: data_buf = 8'h43;
			13'h0d72: data_buf = 8'h0d;
			13'h0d73: data_buf = 8'hfe;
			13'h0d74: data_buf = 8'h2e;
			13'h0d75: data_buf = 8'hca;
			13'h0d76: data_buf = 8'ha3;
			13'h0d77: data_buf = 8'h17;
			13'h0d78: data_buf = 8'hfe;
			13'h0d79: data_buf = 8'had;
			13'h0d7a: data_buf = 8'hca;
			13'h0d7b: data_buf = 8'h99;
			13'h0d7c: data_buf = 8'h0d;
			13'h0d7d: data_buf = 8'hfe;
			13'h0d7e: data_buf = 8'h22;
			13'h0d7f: data_buf = 8'hca;
			13'h0d80: data_buf = 8'h52;
			13'h0d81: data_buf = 8'h11;
			13'h0d82: data_buf = 8'hfe;
			13'h0d83: data_buf = 8'haa;
			13'h0d84: data_buf = 8'hca;
			13'h0d85: data_buf = 8'h8b;
			13'h0d86: data_buf = 8'h0e;
			13'h0d87: data_buf = 8'hfe;
			13'h0d88: data_buf = 8'ha7;
			13'h0d89: data_buf = 8'hca;
			13'h0d8a: data_buf = 8'hb6;
			13'h0d8b: data_buf = 8'h10;
			13'h0d8c: data_buf = 8'hd6;
			13'h0d8d: data_buf = 8'hb6;
			13'h0d8e: data_buf = 8'hd2;
			13'h0d8f: data_buf = 8'hbb;
			13'h0d90: data_buf = 8'h0d;
			13'h0d91: data_buf = 8'hcd;
			13'h0d92: data_buf = 8'hc8;
			13'h0d93: data_buf = 8'h0c;
			13'h0d94: data_buf = 8'hcd;
			13'h0d95: data_buf = 8'hc3;
			13'h0d96: data_buf = 8'h06;
			13'h0d97: data_buf = 8'h29;
			13'h0d98: data_buf = 8'hc9;
			13'h0d99: data_buf = 8'h16;
			13'h0d9a: data_buf = 8'h7d;
			13'h0d9b: data_buf = 8'hcd;
			13'h0d9c: data_buf = 8'hcf;
			13'h0d9d: data_buf = 8'h0c;
			13'h0d9e: data_buf = 8'h2a;
			13'h0d9f: data_buf = 8'h15;
			13'h0da0: data_buf = 8'h81;
			13'h0da1: data_buf = 8'he5;
			13'h0da2: data_buf = 8'hcd;
			13'h0da3: data_buf = 8'hc5;
			13'h0da4: data_buf = 8'h16;
			13'h0da5: data_buf = 8'hcd;
			13'h0da6: data_buf = 8'hbd;
			13'h0da7: data_buf = 8'h0c;
			13'h0da8: data_buf = 8'he1;
			13'h0da9: data_buf = 8'hc9;
			13'h0daa: data_buf = 8'hcd;
			13'h0dab: data_buf = 8'hb0;
			13'h0dac: data_buf = 8'h0e;
			13'h0dad: data_buf = 8'he5;
			13'h0dae: data_buf = 8'heb;
			13'h0daf: data_buf = 8'h22;
			13'h0db0: data_buf = 8'h29;
			13'h0db1: data_buf = 8'h81;
			13'h0db2: data_buf = 8'h3a;
			13'h0db3: data_buf = 8'hf2;
			13'h0db4: data_buf = 8'h80;
			13'h0db5: data_buf = 8'hb7;
			13'h0db6: data_buf = 8'hcc;
			13'h0db7: data_buf = 8'hda;
			13'h0db8: data_buf = 8'h16;
			13'h0db9: data_buf = 8'he1;
			13'h0dba: data_buf = 8'hc9;
			13'h0dbb: data_buf = 8'h06;
			13'h0dbc: data_buf = 8'h00;
			13'h0dbd: data_buf = 8'h07;
			13'h0dbe: data_buf = 8'h4f;
			13'h0dbf: data_buf = 8'hc5;
			13'h0dc0: data_buf = 8'hcd;
			13'h0dc1: data_buf = 8'h4d;
			13'h0dc2: data_buf = 8'h08;
			13'h0dc3: data_buf = 8'h79;
			13'h0dc4: data_buf = 8'hfe;
			13'h0dc5: data_buf = 8'h31;
			13'h0dc6: data_buf = 8'hda;
			13'h0dc7: data_buf = 8'he2;
			13'h0dc8: data_buf = 8'h0d;
			13'h0dc9: data_buf = 8'hcd;
			13'h0dca: data_buf = 8'hc8;
			13'h0dcb: data_buf = 8'h0c;
			13'h0dcc: data_buf = 8'hcd;
			13'h0dcd: data_buf = 8'hc3;
			13'h0dce: data_buf = 8'h06;
			13'h0dcf: data_buf = 8'h2c;
			13'h0dd0: data_buf = 8'hcd;
			13'h0dd1: data_buf = 8'hbe;
			13'h0dd2: data_buf = 8'h0c;
			13'h0dd3: data_buf = 8'heb;
			13'h0dd4: data_buf = 8'h2a;
			13'h0dd5: data_buf = 8'h29;
			13'h0dd6: data_buf = 8'h81;
			13'h0dd7: data_buf = 8'he3;
			13'h0dd8: data_buf = 8'he5;
			13'h0dd9: data_buf = 8'heb;
			13'h0dda: data_buf = 8'hcd;
			13'h0ddb: data_buf = 8'h1b;
			13'h0ddc: data_buf = 8'h14;
			13'h0ddd: data_buf = 8'heb;
			13'h0dde: data_buf = 8'he3;
			13'h0ddf: data_buf = 8'hc3;
			13'h0de0: data_buf = 8'hea;
			13'h0de1: data_buf = 8'h0d;
			13'h0de2: data_buf = 8'hcd;
			13'h0de3: data_buf = 8'h91;
			13'h0de4: data_buf = 8'h0d;
			13'h0de5: data_buf = 8'he3;
			13'h0de6: data_buf = 8'h11;
			13'h0de7: data_buf = 8'ha5;
			13'h0de8: data_buf = 8'h0d;
			13'h0de9: data_buf = 8'hd5;
			13'h0dea: data_buf = 8'h01;
			13'h0deb: data_buf = 8'h46;
			13'h0dec: data_buf = 8'h01;
			13'h0ded: data_buf = 8'h09;
			13'h0dee: data_buf = 8'h4e;
			13'h0def: data_buf = 8'h23;
			13'h0df0: data_buf = 8'h66;
			13'h0df1: data_buf = 8'h69;
			13'h0df2: data_buf = 8'he9;
			13'h0df3: data_buf = 8'h15;
			13'h0df4: data_buf = 8'hfe;
			13'h0df5: data_buf = 8'had;
			13'h0df6: data_buf = 8'hc8;
			13'h0df7: data_buf = 8'hfe;
			13'h0df8: data_buf = 8'h2d;
			13'h0df9: data_buf = 8'hc8;
			13'h0dfa: data_buf = 8'h14;
			13'h0dfb: data_buf = 8'hfe;
			13'h0dfc: data_buf = 8'h2b;
			13'h0dfd: data_buf = 8'hc8;
			13'h0dfe: data_buf = 8'hfe;
			13'h0dff: data_buf = 8'hac;
			13'h0e00: data_buf = 8'hc8;
			13'h0e01: data_buf = 8'h2b;
			13'h0e02: data_buf = 8'hc9;
			13'h0e03: data_buf = 8'hf6;
			13'h0e04: data_buf = 8'haf;
			13'h0e05: data_buf = 8'hf5;
			13'h0e06: data_buf = 8'hcd;
			13'h0e07: data_buf = 8'hbd;
			13'h0e08: data_buf = 8'h0c;
			13'h0e09: data_buf = 8'hcd;
			13'h0e0a: data_buf = 8'hff;
			13'h0e0b: data_buf = 8'h08;
			13'h0e0c: data_buf = 8'hf1;
			13'h0e0d: data_buf = 8'heb;
			13'h0e0e: data_buf = 8'hc1;
			13'h0e0f: data_buf = 8'he3;
			13'h0e10: data_buf = 8'heb;
			13'h0e11: data_buf = 8'hcd;
			13'h0e12: data_buf = 8'hdd;
			13'h0e13: data_buf = 8'h16;
			13'h0e14: data_buf = 8'hf5;
			13'h0e15: data_buf = 8'hcd;
			13'h0e16: data_buf = 8'hff;
			13'h0e17: data_buf = 8'h08;
			13'h0e18: data_buf = 8'hf1;
			13'h0e19: data_buf = 8'hc1;
			13'h0e1a: data_buf = 8'h79;
			13'h0e1b: data_buf = 8'h21;
			13'h0e1c: data_buf = 8'h74;
			13'h0e1d: data_buf = 8'h10;
			13'h0e1e: data_buf = 8'hc2;
			13'h0e1f: data_buf = 8'h26;
			13'h0e20: data_buf = 8'h0e;
			13'h0e21: data_buf = 8'ha3;
			13'h0e22: data_buf = 8'h4f;
			13'h0e23: data_buf = 8'h78;
			13'h0e24: data_buf = 8'ha2;
			13'h0e25: data_buf = 8'he9;
			13'h0e26: data_buf = 8'hb3;
			13'h0e27: data_buf = 8'h4f;
			13'h0e28: data_buf = 8'h78;
			13'h0e29: data_buf = 8'hb2;
			13'h0e2a: data_buf = 8'he9;
			13'h0e2b: data_buf = 8'h21;
			13'h0e2c: data_buf = 8'h3d;
			13'h0e2d: data_buf = 8'h0e;
			13'h0e2e: data_buf = 8'h3a;
			13'h0e2f: data_buf = 8'hf2;
			13'h0e30: data_buf = 8'h80;
			13'h0e31: data_buf = 8'h1f;
			13'h0e32: data_buf = 8'h7a;
			13'h0e33: data_buf = 8'h17;
			13'h0e34: data_buf = 8'h5f;
			13'h0e35: data_buf = 8'h16;
			13'h0e36: data_buf = 8'h64;
			13'h0e37: data_buf = 8'h78;
			13'h0e38: data_buf = 8'hba;
			13'h0e39: data_buf = 8'hd0;
			13'h0e3a: data_buf = 8'hc3;
			13'h0e3b: data_buf = 8'h2c;
			13'h0e3c: data_buf = 8'h0d;
			13'h0e3d: data_buf = 8'h3f;
			13'h0e3e: data_buf = 8'h0e;
			13'h0e3f: data_buf = 8'h79;
			13'h0e40: data_buf = 8'hb7;
			13'h0e41: data_buf = 8'h1f;
			13'h0e42: data_buf = 8'hc1;
			13'h0e43: data_buf = 8'hd1;
			13'h0e44: data_buf = 8'hf5;
			13'h0e45: data_buf = 8'hcd;
			13'h0e46: data_buf = 8'hbf;
			13'h0e47: data_buf = 8'h0c;
			13'h0e48: data_buf = 8'h21;
			13'h0e49: data_buf = 8'h81;
			13'h0e4a: data_buf = 8'h0e;
			13'h0e4b: data_buf = 8'he5;
			13'h0e4c: data_buf = 8'hca;
			13'h0e4d: data_buf = 8'h17;
			13'h0e4e: data_buf = 8'h17;
			13'h0e4f: data_buf = 8'haf;
			13'h0e50: data_buf = 8'h32;
			13'h0e51: data_buf = 8'hf2;
			13'h0e52: data_buf = 8'h80;
			13'h0e53: data_buf = 8'hd5;
			13'h0e54: data_buf = 8'hcd;
			13'h0e55: data_buf = 8'hd6;
			13'h0e56: data_buf = 8'h12;
			13'h0e57: data_buf = 8'h7e;
			13'h0e58: data_buf = 8'h23;
			13'h0e59: data_buf = 8'h23;
			13'h0e5a: data_buf = 8'h4e;
			13'h0e5b: data_buf = 8'h23;
			13'h0e5c: data_buf = 8'h46;
			13'h0e5d: data_buf = 8'hd1;
			13'h0e5e: data_buf = 8'hc5;
			13'h0e5f: data_buf = 8'hf5;
			13'h0e60: data_buf = 8'hcd;
			13'h0e61: data_buf = 8'hda;
			13'h0e62: data_buf = 8'h12;
			13'h0e63: data_buf = 8'hcd;
			13'h0e64: data_buf = 8'heb;
			13'h0e65: data_buf = 8'h16;
			13'h0e66: data_buf = 8'hf1;
			13'h0e67: data_buf = 8'h57;
			13'h0e68: data_buf = 8'he1;
			13'h0e69: data_buf = 8'h7b;
			13'h0e6a: data_buf = 8'hb2;
			13'h0e6b: data_buf = 8'hc8;
			13'h0e6c: data_buf = 8'h7a;
			13'h0e6d: data_buf = 8'hd6;
			13'h0e6e: data_buf = 8'h01;
			13'h0e6f: data_buf = 8'hd8;
			13'h0e70: data_buf = 8'haf;
			13'h0e71: data_buf = 8'hbb;
			13'h0e72: data_buf = 8'h3c;
			13'h0e73: data_buf = 8'hd0;
			13'h0e74: data_buf = 8'h15;
			13'h0e75: data_buf = 8'h1d;
			13'h0e76: data_buf = 8'h0a;
			13'h0e77: data_buf = 8'hbe;
			13'h0e78: data_buf = 8'h23;
			13'h0e79: data_buf = 8'h03;
			13'h0e7a: data_buf = 8'hca;
			13'h0e7b: data_buf = 8'h69;
			13'h0e7c: data_buf = 8'h0e;
			13'h0e7d: data_buf = 8'h3f;
			13'h0e7e: data_buf = 8'hc3;
			13'h0e7f: data_buf = 8'ha7;
			13'h0e80: data_buf = 8'h16;
			13'h0e81: data_buf = 8'h3c;
			13'h0e82: data_buf = 8'h8f;
			13'h0e83: data_buf = 8'hc1;
			13'h0e84: data_buf = 8'ha0;
			13'h0e85: data_buf = 8'hc6;
			13'h0e86: data_buf = 8'hff;
			13'h0e87: data_buf = 8'h9f;
			13'h0e88: data_buf = 8'hc3;
			13'h0e89: data_buf = 8'hae;
			13'h0e8a: data_buf = 8'h16;
			13'h0e8b: data_buf = 8'h16;
			13'h0e8c: data_buf = 8'h5a;
			13'h0e8d: data_buf = 8'hcd;
			13'h0e8e: data_buf = 8'hcf;
			13'h0e8f: data_buf = 8'h0c;
			13'h0e90: data_buf = 8'hcd;
			13'h0e91: data_buf = 8'hbd;
			13'h0e92: data_buf = 8'h0c;
			13'h0e93: data_buf = 8'hcd;
			13'h0e94: data_buf = 8'hff;
			13'h0e95: data_buf = 8'h08;
			13'h0e96: data_buf = 8'h7b;
			13'h0e97: data_buf = 8'h2f;
			13'h0e98: data_buf = 8'h4f;
			13'h0e99: data_buf = 8'h7a;
			13'h0e9a: data_buf = 8'h2f;
			13'h0e9b: data_buf = 8'hcd;
			13'h0e9c: data_buf = 8'h74;
			13'h0e9d: data_buf = 8'h10;
			13'h0e9e: data_buf = 8'hc1;
			13'h0e9f: data_buf = 8'hc3;
			13'h0ea0: data_buf = 8'hdb;
			13'h0ea1: data_buf = 8'h0c;
			13'h0ea2: data_buf = 8'h2b;
			13'h0ea3: data_buf = 8'hcd;
			13'h0ea4: data_buf = 8'h4d;
			13'h0ea5: data_buf = 8'h08;
			13'h0ea6: data_buf = 8'hc8;
			13'h0ea7: data_buf = 8'hcd;
			13'h0ea8: data_buf = 8'hc3;
			13'h0ea9: data_buf = 8'h06;
			13'h0eaa: data_buf = 8'h2c;
			13'h0eab: data_buf = 8'h01;
			13'h0eac: data_buf = 8'ha2;
			13'h0ead: data_buf = 8'h0e;
			13'h0eae: data_buf = 8'hc5;
			13'h0eaf: data_buf = 8'hf6;
			13'h0eb0: data_buf = 8'haf;
			13'h0eb1: data_buf = 8'h32;
			13'h0eb2: data_buf = 8'hf1;
			13'h0eb3: data_buf = 8'h80;
			13'h0eb4: data_buf = 8'h46;
			13'h0eb5: data_buf = 8'hcd;
			13'h0eb6: data_buf = 8'heb;
			13'h0eb7: data_buf = 8'h08;
			13'h0eb8: data_buf = 8'hda;
			13'h0eb9: data_buf = 8'hf5;
			13'h0eba: data_buf = 8'h03;
			13'h0ebb: data_buf = 8'haf;
			13'h0ebc: data_buf = 8'h4f;
			13'h0ebd: data_buf = 8'h32;
			13'h0ebe: data_buf = 8'hf2;
			13'h0ebf: data_buf = 8'h80;
			13'h0ec0: data_buf = 8'hcd;
			13'h0ec1: data_buf = 8'h4d;
			13'h0ec2: data_buf = 8'h08;
			13'h0ec3: data_buf = 8'hda;
			13'h0ec4: data_buf = 8'hcc;
			13'h0ec5: data_buf = 8'h0e;
			13'h0ec6: data_buf = 8'hcd;
			13'h0ec7: data_buf = 8'heb;
			13'h0ec8: data_buf = 8'h08;
			13'h0ec9: data_buf = 8'hda;
			13'h0eca: data_buf = 8'hd9;
			13'h0ecb: data_buf = 8'h0e;
			13'h0ecc: data_buf = 8'h4f;
			13'h0ecd: data_buf = 8'hcd;
			13'h0ece: data_buf = 8'h4d;
			13'h0ecf: data_buf = 8'h08;
			13'h0ed0: data_buf = 8'hda;
			13'h0ed1: data_buf = 8'hcd;
			13'h0ed2: data_buf = 8'h0e;
			13'h0ed3: data_buf = 8'hcd;
			13'h0ed4: data_buf = 8'heb;
			13'h0ed5: data_buf = 8'h08;
			13'h0ed6: data_buf = 8'hd2;
			13'h0ed7: data_buf = 8'hcd;
			13'h0ed8: data_buf = 8'h0e;
			13'h0ed9: data_buf = 8'hd6;
			13'h0eda: data_buf = 8'h24;
			13'h0edb: data_buf = 8'hc2;
			13'h0edc: data_buf = 8'he8;
			13'h0edd: data_buf = 8'h0e;
			13'h0ede: data_buf = 8'h3c;
			13'h0edf: data_buf = 8'h32;
			13'h0ee0: data_buf = 8'hf2;
			13'h0ee1: data_buf = 8'h80;
			13'h0ee2: data_buf = 8'h0f;
			13'h0ee3: data_buf = 8'h81;
			13'h0ee4: data_buf = 8'h4f;
			13'h0ee5: data_buf = 8'hcd;
			13'h0ee6: data_buf = 8'h4d;
			13'h0ee7: data_buf = 8'h08;
			13'h0ee8: data_buf = 8'h3a;
			13'h0ee9: data_buf = 8'h10;
			13'h0eea: data_buf = 8'h81;
			13'h0eeb: data_buf = 8'h3d;
			13'h0eec: data_buf = 8'hca;
			13'h0eed: data_buf = 8'h95;
			13'h0eee: data_buf = 8'h0f;
			13'h0eef: data_buf = 8'hf2;
			13'h0ef0: data_buf = 8'hf8;
			13'h0ef1: data_buf = 8'h0e;
			13'h0ef2: data_buf = 8'h7e;
			13'h0ef3: data_buf = 8'hd6;
			13'h0ef4: data_buf = 8'h28;
			13'h0ef5: data_buf = 8'hca;
			13'h0ef6: data_buf = 8'h6d;
			13'h0ef7: data_buf = 8'h0f;
			13'h0ef8: data_buf = 8'haf;
			13'h0ef9: data_buf = 8'h32;
			13'h0efa: data_buf = 8'h10;
			13'h0efb: data_buf = 8'h81;
			13'h0efc: data_buf = 8'he5;
			13'h0efd: data_buf = 8'h50;
			13'h0efe: data_buf = 8'h59;
			13'h0eff: data_buf = 8'h2a;
			13'h0f00: data_buf = 8'h23;
			13'h0f01: data_buf = 8'h81;
			13'h0f02: data_buf = 8'hcd;
			13'h0f03: data_buf = 8'hbd;
			13'h0f04: data_buf = 8'h06;
			13'h0f05: data_buf = 8'h11;
			13'h0f06: data_buf = 8'h25;
			13'h0f07: data_buf = 8'h81;
			13'h0f08: data_buf = 8'hca;
			13'h0f09: data_buf = 8'hdd;
			13'h0f0a: data_buf = 8'h15;
			13'h0f0b: data_buf = 8'h2a;
			13'h0f0c: data_buf = 8'h1d;
			13'h0f0d: data_buf = 8'h81;
			13'h0f0e: data_buf = 8'heb;
			13'h0f0f: data_buf = 8'h2a;
			13'h0f10: data_buf = 8'h1b;
			13'h0f11: data_buf = 8'h81;
			13'h0f12: data_buf = 8'hcd;
			13'h0f13: data_buf = 8'hbd;
			13'h0f14: data_buf = 8'h06;
			13'h0f15: data_buf = 8'hca;
			13'h0f16: data_buf = 8'h2b;
			13'h0f17: data_buf = 8'h0f;
			13'h0f18: data_buf = 8'h79;
			13'h0f19: data_buf = 8'h96;
			13'h0f1a: data_buf = 8'h23;
			13'h0f1b: data_buf = 8'hc2;
			13'h0f1c: data_buf = 8'h20;
			13'h0f1d: data_buf = 8'h0f;
			13'h0f1e: data_buf = 8'h78;
			13'h0f1f: data_buf = 8'h96;
			13'h0f20: data_buf = 8'h23;
			13'h0f21: data_buf = 8'hca;
			13'h0f22: data_buf = 8'h5f;
			13'h0f23: data_buf = 8'h0f;
			13'h0f24: data_buf = 8'h23;
			13'h0f25: data_buf = 8'h23;
			13'h0f26: data_buf = 8'h23;
			13'h0f27: data_buf = 8'h23;
			13'h0f28: data_buf = 8'hc3;
			13'h0f29: data_buf = 8'h12;
			13'h0f2a: data_buf = 8'h0f;
			13'h0f2b: data_buf = 8'he1;
			13'h0f2c: data_buf = 8'he3;
			13'h0f2d: data_buf = 8'hd5;
			13'h0f2e: data_buf = 8'h11;
			13'h0f2f: data_buf = 8'had;
			13'h0f30: data_buf = 8'h0d;
			13'h0f31: data_buf = 8'hcd;
			13'h0f32: data_buf = 8'hbd;
			13'h0f33: data_buf = 8'h06;
			13'h0f34: data_buf = 8'hd1;
			13'h0f35: data_buf = 8'hca;
			13'h0f36: data_buf = 8'h62;
			13'h0f37: data_buf = 8'h0f;
			13'h0f38: data_buf = 8'he3;
			13'h0f39: data_buf = 8'he5;
			13'h0f3a: data_buf = 8'hc5;
			13'h0f3b: data_buf = 8'h01;
			13'h0f3c: data_buf = 8'h06;
			13'h0f3d: data_buf = 8'h00;
			13'h0f3e: data_buf = 8'h2a;
			13'h0f3f: data_buf = 8'h1f;
			13'h0f40: data_buf = 8'h81;
			13'h0f41: data_buf = 8'he5;
			13'h0f42: data_buf = 8'h09;
			13'h0f43: data_buf = 8'hc1;
			13'h0f44: data_buf = 8'he5;
			13'h0f45: data_buf = 8'hcd;
			13'h0f46: data_buf = 8'hc1;
			13'h0f47: data_buf = 8'h03;
			13'h0f48: data_buf = 8'he1;
			13'h0f49: data_buf = 8'h22;
			13'h0f4a: data_buf = 8'h1f;
			13'h0f4b: data_buf = 8'h81;
			13'h0f4c: data_buf = 8'h60;
			13'h0f4d: data_buf = 8'h69;
			13'h0f4e: data_buf = 8'h22;
			13'h0f4f: data_buf = 8'h1d;
			13'h0f50: data_buf = 8'h81;
			13'h0f51: data_buf = 8'h2b;
			13'h0f52: data_buf = 8'h36;
			13'h0f53: data_buf = 8'h00;
			13'h0f54: data_buf = 8'hcd;
			13'h0f55: data_buf = 8'hbd;
			13'h0f56: data_buf = 8'h06;
			13'h0f57: data_buf = 8'hc2;
			13'h0f58: data_buf = 8'h51;
			13'h0f59: data_buf = 8'h0f;
			13'h0f5a: data_buf = 8'hd1;
			13'h0f5b: data_buf = 8'h73;
			13'h0f5c: data_buf = 8'h23;
			13'h0f5d: data_buf = 8'h72;
			13'h0f5e: data_buf = 8'h23;
			13'h0f5f: data_buf = 8'heb;
			13'h0f60: data_buf = 8'he1;
			13'h0f61: data_buf = 8'hc9;
			13'h0f62: data_buf = 8'h32;
			13'h0f63: data_buf = 8'h2c;
			13'h0f64: data_buf = 8'h81;
			13'h0f65: data_buf = 8'h21;
			13'h0f66: data_buf = 8'h91;
			13'h0f67: data_buf = 8'h03;
			13'h0f68: data_buf = 8'h22;
			13'h0f69: data_buf = 8'h29;
			13'h0f6a: data_buf = 8'h81;
			13'h0f6b: data_buf = 8'he1;
			13'h0f6c: data_buf = 8'hc9;
			13'h0f6d: data_buf = 8'he5;
			13'h0f6e: data_buf = 8'h2a;
			13'h0f6f: data_buf = 8'hf1;
			13'h0f70: data_buf = 8'h80;
			13'h0f71: data_buf = 8'he3;
			13'h0f72: data_buf = 8'h57;
			13'h0f73: data_buf = 8'hd5;
			13'h0f74: data_buf = 8'hc5;
			13'h0f75: data_buf = 8'hcd;
			13'h0f76: data_buf = 8'hf3;
			13'h0f77: data_buf = 8'h08;
			13'h0f78: data_buf = 8'hc1;
			13'h0f79: data_buf = 8'hf1;
			13'h0f7a: data_buf = 8'heb;
			13'h0f7b: data_buf = 8'he3;
			13'h0f7c: data_buf = 8'he5;
			13'h0f7d: data_buf = 8'heb;
			13'h0f7e: data_buf = 8'h3c;
			13'h0f7f: data_buf = 8'h57;
			13'h0f80: data_buf = 8'h7e;
			13'h0f81: data_buf = 8'hfe;
			13'h0f82: data_buf = 8'h2c;
			13'h0f83: data_buf = 8'hca;
			13'h0f84: data_buf = 8'h73;
			13'h0f85: data_buf = 8'h0f;
			13'h0f86: data_buf = 8'hcd;
			13'h0f87: data_buf = 8'hc3;
			13'h0f88: data_buf = 8'h06;
			13'h0f89: data_buf = 8'h29;
			13'h0f8a: data_buf = 8'h22;
			13'h0f8b: data_buf = 8'h15;
			13'h0f8c: data_buf = 8'h81;
			13'h0f8d: data_buf = 8'he1;
			13'h0f8e: data_buf = 8'h22;
			13'h0f8f: data_buf = 8'hf1;
			13'h0f90: data_buf = 8'h80;
			13'h0f91: data_buf = 8'h1e;
			13'h0f92: data_buf = 8'h00;
			13'h0f93: data_buf = 8'hd5;
			13'h0f94: data_buf = 8'h11;
			13'h0f95: data_buf = 8'he5;
			13'h0f96: data_buf = 8'hf5;
			13'h0f97: data_buf = 8'h2a;
			13'h0f98: data_buf = 8'h1d;
			13'h0f99: data_buf = 8'h81;
			13'h0f9a: data_buf = 8'h3e;
			13'h0f9b: data_buf = 8'h19;
			13'h0f9c: data_buf = 8'heb;
			13'h0f9d: data_buf = 8'h2a;
			13'h0f9e: data_buf = 8'h1f;
			13'h0f9f: data_buf = 8'h81;
			13'h0fa0: data_buf = 8'heb;
			13'h0fa1: data_buf = 8'hcd;
			13'h0fa2: data_buf = 8'hbd;
			13'h0fa3: data_buf = 8'h06;
			13'h0fa4: data_buf = 8'hca;
			13'h0fa5: data_buf = 8'hcd;
			13'h0fa6: data_buf = 8'h0f;
			13'h0fa7: data_buf = 8'h7e;
			13'h0fa8: data_buf = 8'hb9;
			13'h0fa9: data_buf = 8'h23;
			13'h0faa: data_buf = 8'hc2;
			13'h0fab: data_buf = 8'haf;
			13'h0fac: data_buf = 8'h0f;
			13'h0fad: data_buf = 8'h7e;
			13'h0fae: data_buf = 8'hb8;
			13'h0faf: data_buf = 8'h23;
			13'h0fb0: data_buf = 8'h5e;
			13'h0fb1: data_buf = 8'h23;
			13'h0fb2: data_buf = 8'h56;
			13'h0fb3: data_buf = 8'h23;
			13'h0fb4: data_buf = 8'hc2;
			13'h0fb5: data_buf = 8'h9b;
			13'h0fb6: data_buf = 8'h0f;
			13'h0fb7: data_buf = 8'h3a;
			13'h0fb8: data_buf = 8'hf1;
			13'h0fb9: data_buf = 8'h80;
			13'h0fba: data_buf = 8'hb7;
			13'h0fbb: data_buf = 8'hc2;
			13'h0fbc: data_buf = 8'hfe;
			13'h0fbd: data_buf = 8'h03;
			13'h0fbe: data_buf = 8'hf1;
			13'h0fbf: data_buf = 8'h44;
			13'h0fc0: data_buf = 8'h4d;
			13'h0fc1: data_buf = 8'hca;
			13'h0fc2: data_buf = 8'hdd;
			13'h0fc3: data_buf = 8'h15;
			13'h0fc4: data_buf = 8'h96;
			13'h0fc5: data_buf = 8'hca;
			13'h0fc6: data_buf = 8'h2b;
			13'h0fc7: data_buf = 8'h10;
			13'h0fc8: data_buf = 8'h1e;
			13'h0fc9: data_buf = 8'h10;
			13'h0fca: data_buf = 8'hc3;
			13'h0fcb: data_buf = 8'h09;
			13'h0fcc: data_buf = 8'h04;
			13'h0fcd: data_buf = 8'h11;
			13'h0fce: data_buf = 8'h04;
			13'h0fcf: data_buf = 8'h00;
			13'h0fd0: data_buf = 8'hf1;
			13'h0fd1: data_buf = 8'hca;
			13'h0fd2: data_buf = 8'h14;
			13'h0fd3: data_buf = 8'h09;
			13'h0fd4: data_buf = 8'h71;
			13'h0fd5: data_buf = 8'h23;
			13'h0fd6: data_buf = 8'h70;
			13'h0fd7: data_buf = 8'h23;
			13'h0fd8: data_buf = 8'h4f;
			13'h0fd9: data_buf = 8'hcd;
			13'h0fda: data_buf = 8'hd2;
			13'h0fdb: data_buf = 8'h03;
			13'h0fdc: data_buf = 8'h23;
			13'h0fdd: data_buf = 8'h23;
			13'h0fde: data_buf = 8'h22;
			13'h0fdf: data_buf = 8'h0a;
			13'h0fe0: data_buf = 8'h81;
			13'h0fe1: data_buf = 8'h71;
			13'h0fe2: data_buf = 8'h23;
			13'h0fe3: data_buf = 8'h3a;
			13'h0fe4: data_buf = 8'hf1;
			13'h0fe5: data_buf = 8'h80;
			13'h0fe6: data_buf = 8'h17;
			13'h0fe7: data_buf = 8'h79;
			13'h0fe8: data_buf = 8'h01;
			13'h0fe9: data_buf = 8'h0b;
			13'h0fea: data_buf = 8'h00;
			13'h0feb: data_buf = 8'hd2;
			13'h0fec: data_buf = 8'hf0;
			13'h0fed: data_buf = 8'h0f;
			13'h0fee: data_buf = 8'hc1;
			13'h0fef: data_buf = 8'h03;
			13'h0ff0: data_buf = 8'h71;
			13'h0ff1: data_buf = 8'h23;
			13'h0ff2: data_buf = 8'h70;
			13'h0ff3: data_buf = 8'h23;
			13'h0ff4: data_buf = 8'hf5;
			13'h0ff5: data_buf = 8'he5;
			13'h0ff6: data_buf = 8'hcd;
			13'h0ff7: data_buf = 8'h88;
			13'h0ff8: data_buf = 8'h17;
			13'h0ff9: data_buf = 8'heb;
			13'h0ffa: data_buf = 8'he1;
			13'h0ffb: data_buf = 8'hf1;
			13'h0ffc: data_buf = 8'h3d;
			13'h0ffd: data_buf = 8'hc2;
			13'h0ffe: data_buf = 8'he8;
			13'h0fff: data_buf = 8'h0f;
			13'h1000: data_buf = 8'hf5;
			13'h1001: data_buf = 8'h42;
			13'h1002: data_buf = 8'h4b;
			13'h1003: data_buf = 8'heb;
			13'h1004: data_buf = 8'h19;
			13'h1005: data_buf = 8'hda;
			13'h1006: data_buf = 8'hea;
			13'h1007: data_buf = 8'h03;
			13'h1008: data_buf = 8'hcd;
			13'h1009: data_buf = 8'hdb;
			13'h100a: data_buf = 8'h03;
			13'h100b: data_buf = 8'h22;
			13'h100c: data_buf = 8'h1f;
			13'h100d: data_buf = 8'h81;
			13'h100e: data_buf = 8'h2b;
			13'h100f: data_buf = 8'h36;
			13'h1010: data_buf = 8'h00;
			13'h1011: data_buf = 8'hcd;
			13'h1012: data_buf = 8'hbd;
			13'h1013: data_buf = 8'h06;
			13'h1014: data_buf = 8'hc2;
			13'h1015: data_buf = 8'h0e;
			13'h1016: data_buf = 8'h10;
			13'h1017: data_buf = 8'h03;
			13'h1018: data_buf = 8'h57;
			13'h1019: data_buf = 8'h2a;
			13'h101a: data_buf = 8'h0a;
			13'h101b: data_buf = 8'h81;
			13'h101c: data_buf = 8'h5e;
			13'h101d: data_buf = 8'heb;
			13'h101e: data_buf = 8'h29;
			13'h101f: data_buf = 8'h09;
			13'h1020: data_buf = 8'heb;
			13'h1021: data_buf = 8'h2b;
			13'h1022: data_buf = 8'h2b;
			13'h1023: data_buf = 8'h73;
			13'h1024: data_buf = 8'h23;
			13'h1025: data_buf = 8'h72;
			13'h1026: data_buf = 8'h23;
			13'h1027: data_buf = 8'hf1;
			13'h1028: data_buf = 8'hda;
			13'h1029: data_buf = 8'h4f;
			13'h102a: data_buf = 8'h10;
			13'h102b: data_buf = 8'h47;
			13'h102c: data_buf = 8'h4f;
			13'h102d: data_buf = 8'h7e;
			13'h102e: data_buf = 8'h23;
			13'h102f: data_buf = 8'h16;
			13'h1030: data_buf = 8'he1;
			13'h1031: data_buf = 8'h5e;
			13'h1032: data_buf = 8'h23;
			13'h1033: data_buf = 8'h56;
			13'h1034: data_buf = 8'h23;
			13'h1035: data_buf = 8'he3;
			13'h1036: data_buf = 8'hf5;
			13'h1037: data_buf = 8'hcd;
			13'h1038: data_buf = 8'hbd;
			13'h1039: data_buf = 8'h06;
			13'h103a: data_buf = 8'hd2;
			13'h103b: data_buf = 8'hc8;
			13'h103c: data_buf = 8'h0f;
			13'h103d: data_buf = 8'he5;
			13'h103e: data_buf = 8'hcd;
			13'h103f: data_buf = 8'h88;
			13'h1040: data_buf = 8'h17;
			13'h1041: data_buf = 8'hd1;
			13'h1042: data_buf = 8'h19;
			13'h1043: data_buf = 8'hf1;
			13'h1044: data_buf = 8'h3d;
			13'h1045: data_buf = 8'h44;
			13'h1046: data_buf = 8'h4d;
			13'h1047: data_buf = 8'hc2;
			13'h1048: data_buf = 8'h30;
			13'h1049: data_buf = 8'h10;
			13'h104a: data_buf = 8'h29;
			13'h104b: data_buf = 8'h29;
			13'h104c: data_buf = 8'hc1;
			13'h104d: data_buf = 8'h09;
			13'h104e: data_buf = 8'heb;
			13'h104f: data_buf = 8'h2a;
			13'h1050: data_buf = 8'h15;
			13'h1051: data_buf = 8'h81;
			13'h1052: data_buf = 8'hc9;
			13'h1053: data_buf = 8'h2a;
			13'h1054: data_buf = 8'h1f;
			13'h1055: data_buf = 8'h81;
			13'h1056: data_buf = 8'heb;
			13'h1057: data_buf = 8'h21;
			13'h1058: data_buf = 8'h00;
			13'h1059: data_buf = 8'h00;
			13'h105a: data_buf = 8'h39;
			13'h105b: data_buf = 8'h3a;
			13'h105c: data_buf = 8'hf2;
			13'h105d: data_buf = 8'h80;
			13'h105e: data_buf = 8'hb7;
			13'h105f: data_buf = 8'hca;
			13'h1060: data_buf = 8'h6f;
			13'h1061: data_buf = 8'h10;
			13'h1062: data_buf = 8'hcd;
			13'h1063: data_buf = 8'hd6;
			13'h1064: data_buf = 8'h12;
			13'h1065: data_buf = 8'hcd;
			13'h1066: data_buf = 8'hd6;
			13'h1067: data_buf = 8'h11;
			13'h1068: data_buf = 8'h2a;
			13'h1069: data_buf = 8'h9f;
			13'h106a: data_buf = 8'h80;
			13'h106b: data_buf = 8'heb;
			13'h106c: data_buf = 8'h2a;
			13'h106d: data_buf = 8'h08;
			13'h106e: data_buf = 8'h81;
			13'h106f: data_buf = 8'h7d;
			13'h1070: data_buf = 8'h93;
			13'h1071: data_buf = 8'h4f;
			13'h1072: data_buf = 8'h7c;
			13'h1073: data_buf = 8'h9a;
			13'h1074: data_buf = 8'h41;
			13'h1075: data_buf = 8'h50;
			13'h1076: data_buf = 8'h1e;
			13'h1077: data_buf = 8'h00;
			13'h1078: data_buf = 8'h21;
			13'h1079: data_buf = 8'hf2;
			13'h107a: data_buf = 8'h80;
			13'h107b: data_buf = 8'h73;
			13'h107c: data_buf = 8'h06;
			13'h107d: data_buf = 8'h90;
			13'h107e: data_buf = 8'hc3;
			13'h107f: data_buf = 8'hb3;
			13'h1080: data_buf = 8'h16;
			13'h1081: data_buf = 8'h3a;
			13'h1082: data_buf = 8'hf0;
			13'h1083: data_buf = 8'h80;
			13'h1084: data_buf = 8'h47;
			13'h1085: data_buf = 8'haf;
			13'h1086: data_buf = 8'hc3;
			13'h1087: data_buf = 8'h75;
			13'h1088: data_buf = 8'h10;
			13'h1089: data_buf = 8'hcd;
			13'h108a: data_buf = 8'h0c;
			13'h108b: data_buf = 8'h11;
			13'h108c: data_buf = 8'hcd;
			13'h108d: data_buf = 8'hfe;
			13'h108e: data_buf = 8'h10;
			13'h108f: data_buf = 8'h01;
			13'h1090: data_buf = 8'he4;
			13'h1091: data_buf = 8'h09;
			13'h1092: data_buf = 8'hc5;
			13'h1093: data_buf = 8'hd5;
			13'h1094: data_buf = 8'hcd;
			13'h1095: data_buf = 8'hc3;
			13'h1096: data_buf = 8'h06;
			13'h1097: data_buf = 8'h28;
			13'h1098: data_buf = 8'hcd;
			13'h1099: data_buf = 8'hb0;
			13'h109a: data_buf = 8'h0e;
			13'h109b: data_buf = 8'he5;
			13'h109c: data_buf = 8'heb;
			13'h109d: data_buf = 8'h2b;
			13'h109e: data_buf = 8'h56;
			13'h109f: data_buf = 8'h2b;
			13'h10a0: data_buf = 8'h5e;
			13'h10a1: data_buf = 8'he1;
			13'h10a2: data_buf = 8'hcd;
			13'h10a3: data_buf = 8'hbd;
			13'h10a4: data_buf = 8'h0c;
			13'h10a5: data_buf = 8'hcd;
			13'h10a6: data_buf = 8'hc3;
			13'h10a7: data_buf = 8'h06;
			13'h10a8: data_buf = 8'h29;
			13'h10a9: data_buf = 8'hcd;
			13'h10aa: data_buf = 8'hc3;
			13'h10ab: data_buf = 8'h06;
			13'h10ac: data_buf = 8'hb4;
			13'h10ad: data_buf = 8'h44;
			13'h10ae: data_buf = 8'h4d;
			13'h10af: data_buf = 8'he3;
			13'h10b0: data_buf = 8'h71;
			13'h10b1: data_buf = 8'h23;
			13'h10b2: data_buf = 8'h70;
			13'h10b3: data_buf = 8'hc3;
			13'h10b4: data_buf = 8'h4b;
			13'h10b5: data_buf = 8'h11;
			13'h10b6: data_buf = 8'hcd;
			13'h10b7: data_buf = 8'h0c;
			13'h10b8: data_buf = 8'h11;
			13'h10b9: data_buf = 8'hd5;
			13'h10ba: data_buf = 8'hcd;
			13'h10bb: data_buf = 8'h91;
			13'h10bc: data_buf = 8'h0d;
			13'h10bd: data_buf = 8'hcd;
			13'h10be: data_buf = 8'hbd;
			13'h10bf: data_buf = 8'h0c;
			13'h10c0: data_buf = 8'he3;
			13'h10c1: data_buf = 8'h5e;
			13'h10c2: data_buf = 8'h23;
			13'h10c3: data_buf = 8'h56;
			13'h10c4: data_buf = 8'h23;
			13'h10c5: data_buf = 8'h7a;
			13'h10c6: data_buf = 8'hb3;
			13'h10c7: data_buf = 8'hca;
			13'h10c8: data_buf = 8'h01;
			13'h10c9: data_buf = 8'h04;
			13'h10ca: data_buf = 8'h7e;
			13'h10cb: data_buf = 8'h23;
			13'h10cc: data_buf = 8'h66;
			13'h10cd: data_buf = 8'h6f;
			13'h10ce: data_buf = 8'he5;
			13'h10cf: data_buf = 8'h2a;
			13'h10d0: data_buf = 8'h23;
			13'h10d1: data_buf = 8'h81;
			13'h10d2: data_buf = 8'he3;
			13'h10d3: data_buf = 8'h22;
			13'h10d4: data_buf = 8'h23;
			13'h10d5: data_buf = 8'h81;
			13'h10d6: data_buf = 8'h2a;
			13'h10d7: data_buf = 8'h27;
			13'h10d8: data_buf = 8'h81;
			13'h10d9: data_buf = 8'he5;
			13'h10da: data_buf = 8'h2a;
			13'h10db: data_buf = 8'h25;
			13'h10dc: data_buf = 8'h81;
			13'h10dd: data_buf = 8'he5;
			13'h10de: data_buf = 8'h21;
			13'h10df: data_buf = 8'h25;
			13'h10e0: data_buf = 8'h81;
			13'h10e1: data_buf = 8'hd5;
			13'h10e2: data_buf = 8'hcd;
			13'h10e3: data_buf = 8'hf4;
			13'h10e4: data_buf = 8'h16;
			13'h10e5: data_buf = 8'he1;
			13'h10e6: data_buf = 8'hcd;
			13'h10e7: data_buf = 8'hba;
			13'h10e8: data_buf = 8'h0c;
			13'h10e9: data_buf = 8'h2b;
			13'h10ea: data_buf = 8'hcd;
			13'h10eb: data_buf = 8'h4d;
			13'h10ec: data_buf = 8'h08;
			13'h10ed: data_buf = 8'hc2;
			13'h10ee: data_buf = 8'hf5;
			13'h10ef: data_buf = 8'h03;
			13'h10f0: data_buf = 8'he1;
			13'h10f1: data_buf = 8'h22;
			13'h10f2: data_buf = 8'h25;
			13'h10f3: data_buf = 8'h81;
			13'h10f4: data_buf = 8'he1;
			13'h10f5: data_buf = 8'h22;
			13'h10f6: data_buf = 8'h27;
			13'h10f7: data_buf = 8'h81;
			13'h10f8: data_buf = 8'he1;
			13'h10f9: data_buf = 8'h22;
			13'h10fa: data_buf = 8'h23;
			13'h10fb: data_buf = 8'h81;
			13'h10fc: data_buf = 8'he1;
			13'h10fd: data_buf = 8'hc9;
			13'h10fe: data_buf = 8'he5;
			13'h10ff: data_buf = 8'h2a;
			13'h1100: data_buf = 8'ha1;
			13'h1101: data_buf = 8'h80;
			13'h1102: data_buf = 8'h23;
			13'h1103: data_buf = 8'h7c;
			13'h1104: data_buf = 8'hb5;
			13'h1105: data_buf = 8'he1;
			13'h1106: data_buf = 8'hc0;
			13'h1107: data_buf = 8'h1e;
			13'h1108: data_buf = 8'h16;
			13'h1109: data_buf = 8'hc3;
			13'h110a: data_buf = 8'h09;
			13'h110b: data_buf = 8'h04;
			13'h110c: data_buf = 8'hcd;
			13'h110d: data_buf = 8'hc3;
			13'h110e: data_buf = 8'h06;
			13'h110f: data_buf = 8'ha7;
			13'h1110: data_buf = 8'h3e;
			13'h1111: data_buf = 8'h80;
			13'h1112: data_buf = 8'h32;
			13'h1113: data_buf = 8'h10;
			13'h1114: data_buf = 8'h81;
			13'h1115: data_buf = 8'hb6;
			13'h1116: data_buf = 8'h47;
			13'h1117: data_buf = 8'hcd;
			13'h1118: data_buf = 8'hb5;
			13'h1119: data_buf = 8'h0e;
			13'h111a: data_buf = 8'hc3;
			13'h111b: data_buf = 8'hbd;
			13'h111c: data_buf = 8'h0c;
			13'h111d: data_buf = 8'hcd;
			13'h111e: data_buf = 8'hbd;
			13'h111f: data_buf = 8'h0c;
			13'h1120: data_buf = 8'hcd;
			13'h1121: data_buf = 8'h41;
			13'h1122: data_buf = 8'h18;
			13'h1123: data_buf = 8'hcd;
			13'h1124: data_buf = 8'h51;
			13'h1125: data_buf = 8'h11;
			13'h1126: data_buf = 8'hcd;
			13'h1127: data_buf = 8'hd6;
			13'h1128: data_buf = 8'h12;
			13'h1129: data_buf = 8'h01;
			13'h112a: data_buf = 8'h31;
			13'h112b: data_buf = 8'h13;
			13'h112c: data_buf = 8'hc5;
			13'h112d: data_buf = 8'h7e;
			13'h112e: data_buf = 8'h23;
			13'h112f: data_buf = 8'h23;
			13'h1130: data_buf = 8'he5;
			13'h1131: data_buf = 8'hcd;
			13'h1132: data_buf = 8'hac;
			13'h1133: data_buf = 8'h11;
			13'h1134: data_buf = 8'he1;
			13'h1135: data_buf = 8'h4e;
			13'h1136: data_buf = 8'h23;
			13'h1137: data_buf = 8'h46;
			13'h1138: data_buf = 8'hcd;
			13'h1139: data_buf = 8'h45;
			13'h113a: data_buf = 8'h11;
			13'h113b: data_buf = 8'he5;
			13'h113c: data_buf = 8'h6f;
			13'h113d: data_buf = 8'hcd;
			13'h113e: data_buf = 8'hc9;
			13'h113f: data_buf = 8'h12;
			13'h1140: data_buf = 8'hd1;
			13'h1141: data_buf = 8'hc9;
			13'h1142: data_buf = 8'hcd;
			13'h1143: data_buf = 8'hac;
			13'h1144: data_buf = 8'h11;
			13'h1145: data_buf = 8'h21;
			13'h1146: data_buf = 8'h04;
			13'h1147: data_buf = 8'h81;
			13'h1148: data_buf = 8'he5;
			13'h1149: data_buf = 8'h77;
			13'h114a: data_buf = 8'h23;
			13'h114b: data_buf = 8'h23;
			13'h114c: data_buf = 8'h73;
			13'h114d: data_buf = 8'h23;
			13'h114e: data_buf = 8'h72;
			13'h114f: data_buf = 8'he1;
			13'h1150: data_buf = 8'hc9;
			13'h1151: data_buf = 8'h2b;
			13'h1152: data_buf = 8'h06;
			13'h1153: data_buf = 8'h22;
			13'h1154: data_buf = 8'h50;
			13'h1155: data_buf = 8'he5;
			13'h1156: data_buf = 8'h0e;
			13'h1157: data_buf = 8'hff;
			13'h1158: data_buf = 8'h23;
			13'h1159: data_buf = 8'h7e;
			13'h115a: data_buf = 8'h0c;
			13'h115b: data_buf = 8'hb7;
			13'h115c: data_buf = 8'hca;
			13'h115d: data_buf = 8'h67;
			13'h115e: data_buf = 8'h11;
			13'h115f: data_buf = 8'hba;
			13'h1160: data_buf = 8'hca;
			13'h1161: data_buf = 8'h67;
			13'h1162: data_buf = 8'h11;
			13'h1163: data_buf = 8'hb8;
			13'h1164: data_buf = 8'hc2;
			13'h1165: data_buf = 8'h58;
			13'h1166: data_buf = 8'h11;
			13'h1167: data_buf = 8'hfe;
			13'h1168: data_buf = 8'h22;
			13'h1169: data_buf = 8'hcc;
			13'h116a: data_buf = 8'h4d;
			13'h116b: data_buf = 8'h08;
			13'h116c: data_buf = 8'he3;
			13'h116d: data_buf = 8'h23;
			13'h116e: data_buf = 8'heb;
			13'h116f: data_buf = 8'h79;
			13'h1170: data_buf = 8'hcd;
			13'h1171: data_buf = 8'h45;
			13'h1172: data_buf = 8'h11;
			13'h1173: data_buf = 8'h11;
			13'h1174: data_buf = 8'h04;
			13'h1175: data_buf = 8'h81;
			13'h1176: data_buf = 8'h2a;
			13'h1177: data_buf = 8'hf6;
			13'h1178: data_buf = 8'h80;
			13'h1179: data_buf = 8'h22;
			13'h117a: data_buf = 8'h29;
			13'h117b: data_buf = 8'h81;
			13'h117c: data_buf = 8'h3e;
			13'h117d: data_buf = 8'h01;
			13'h117e: data_buf = 8'h32;
			13'h117f: data_buf = 8'hf2;
			13'h1180: data_buf = 8'h80;
			13'h1181: data_buf = 8'hcd;
			13'h1182: data_buf = 8'hf7;
			13'h1183: data_buf = 8'h16;
			13'h1184: data_buf = 8'hcd;
			13'h1185: data_buf = 8'hbd;
			13'h1186: data_buf = 8'h06;
			13'h1187: data_buf = 8'h22;
			13'h1188: data_buf = 8'hf6;
			13'h1189: data_buf = 8'h80;
			13'h118a: data_buf = 8'he1;
			13'h118b: data_buf = 8'h7e;
			13'h118c: data_buf = 8'hc0;
			13'h118d: data_buf = 8'h1e;
			13'h118e: data_buf = 8'h1e;
			13'h118f: data_buf = 8'hc3;
			13'h1190: data_buf = 8'h09;
			13'h1191: data_buf = 8'h04;
			13'h1192: data_buf = 8'h23;
			13'h1193: data_buf = 8'hcd;
			13'h1194: data_buf = 8'h51;
			13'h1195: data_buf = 8'h11;
			13'h1196: data_buf = 8'hcd;
			13'h1197: data_buf = 8'hd6;
			13'h1198: data_buf = 8'h12;
			13'h1199: data_buf = 8'hcd;
			13'h119a: data_buf = 8'heb;
			13'h119b: data_buf = 8'h16;
			13'h119c: data_buf = 8'h1c;
			13'h119d: data_buf = 8'h1d;
			13'h119e: data_buf = 8'hc8;
			13'h119f: data_buf = 8'h0a;
			13'h11a0: data_buf = 8'hcd;
			13'h11a1: data_buf = 8'hce;
			13'h11a2: data_buf = 8'h06;
			13'h11a3: data_buf = 8'hfe;
			13'h11a4: data_buf = 8'h0d;
			13'h11a5: data_buf = 8'hcc;
			13'h11a6: data_buf = 8'hff;
			13'h11a7: data_buf = 8'h0a;
			13'h11a8: data_buf = 8'h03;
			13'h11a9: data_buf = 8'hc3;
			13'h11aa: data_buf = 8'h9d;
			13'h11ab: data_buf = 8'h11;
			13'h11ac: data_buf = 8'hb7;
			13'h11ad: data_buf = 8'h0e;
			13'h11ae: data_buf = 8'hf1;
			13'h11af: data_buf = 8'hf5;
			13'h11b0: data_buf = 8'h2a;
			13'h11b1: data_buf = 8'h9f;
			13'h11b2: data_buf = 8'h80;
			13'h11b3: data_buf = 8'heb;
			13'h11b4: data_buf = 8'h2a;
			13'h11b5: data_buf = 8'h08;
			13'h11b6: data_buf = 8'h81;
			13'h11b7: data_buf = 8'h2f;
			13'h11b8: data_buf = 8'h4f;
			13'h11b9: data_buf = 8'h06;
			13'h11ba: data_buf = 8'hff;
			13'h11bb: data_buf = 8'h09;
			13'h11bc: data_buf = 8'h23;
			13'h11bd: data_buf = 8'hcd;
			13'h11be: data_buf = 8'hbd;
			13'h11bf: data_buf = 8'h06;
			13'h11c0: data_buf = 8'hda;
			13'h11c1: data_buf = 8'hca;
			13'h11c2: data_buf = 8'h11;
			13'h11c3: data_buf = 8'h22;
			13'h11c4: data_buf = 8'h08;
			13'h11c5: data_buf = 8'h81;
			13'h11c6: data_buf = 8'h23;
			13'h11c7: data_buf = 8'heb;
			13'h11c8: data_buf = 8'hf1;
			13'h11c9: data_buf = 8'hc9;
			13'h11ca: data_buf = 8'hf1;
			13'h11cb: data_buf = 8'h1e;
			13'h11cc: data_buf = 8'h1a;
			13'h11cd: data_buf = 8'hca;
			13'h11ce: data_buf = 8'h09;
			13'h11cf: data_buf = 8'h04;
			13'h11d0: data_buf = 8'hbf;
			13'h11d1: data_buf = 8'hf5;
			13'h11d2: data_buf = 8'h01;
			13'h11d3: data_buf = 8'hae;
			13'h11d4: data_buf = 8'h11;
			13'h11d5: data_buf = 8'hc5;
			13'h11d6: data_buf = 8'h2a;
			13'h11d7: data_buf = 8'hf4;
			13'h11d8: data_buf = 8'h80;
			13'h11d9: data_buf = 8'h22;
			13'h11da: data_buf = 8'h08;
			13'h11db: data_buf = 8'h81;
			13'h11dc: data_buf = 8'h21;
			13'h11dd: data_buf = 8'h00;
			13'h11de: data_buf = 8'h00;
			13'h11df: data_buf = 8'he5;
			13'h11e0: data_buf = 8'h2a;
			13'h11e1: data_buf = 8'h9f;
			13'h11e2: data_buf = 8'h80;
			13'h11e3: data_buf = 8'he5;
			13'h11e4: data_buf = 8'h21;
			13'h11e5: data_buf = 8'hf8;
			13'h11e6: data_buf = 8'h80;
			13'h11e7: data_buf = 8'heb;
			13'h11e8: data_buf = 8'h2a;
			13'h11e9: data_buf = 8'hf6;
			13'h11ea: data_buf = 8'h80;
			13'h11eb: data_buf = 8'heb;
			13'h11ec: data_buf = 8'hcd;
			13'h11ed: data_buf = 8'hbd;
			13'h11ee: data_buf = 8'h06;
			13'h11ef: data_buf = 8'h01;
			13'h11f0: data_buf = 8'he7;
			13'h11f1: data_buf = 8'h11;
			13'h11f2: data_buf = 8'hc2;
			13'h11f3: data_buf = 8'h3b;
			13'h11f4: data_buf = 8'h12;
			13'h11f5: data_buf = 8'h2a;
			13'h11f6: data_buf = 8'h1b;
			13'h11f7: data_buf = 8'h81;
			13'h11f8: data_buf = 8'heb;
			13'h11f9: data_buf = 8'h2a;
			13'h11fa: data_buf = 8'h1d;
			13'h11fb: data_buf = 8'h81;
			13'h11fc: data_buf = 8'heb;
			13'h11fd: data_buf = 8'hcd;
			13'h11fe: data_buf = 8'hbd;
			13'h11ff: data_buf = 8'h06;
			13'h1200: data_buf = 8'hca;
			13'h1201: data_buf = 8'h0e;
			13'h1202: data_buf = 8'h12;
			13'h1203: data_buf = 8'h7e;
			13'h1204: data_buf = 8'h23;
			13'h1205: data_buf = 8'h23;
			13'h1206: data_buf = 8'hb7;
			13'h1207: data_buf = 8'hcd;
			13'h1208: data_buf = 8'h3e;
			13'h1209: data_buf = 8'h12;
			13'h120a: data_buf = 8'hc3;
			13'h120b: data_buf = 8'hf8;
			13'h120c: data_buf = 8'h11;
			13'h120d: data_buf = 8'hc1;
			13'h120e: data_buf = 8'heb;
			13'h120f: data_buf = 8'h2a;
			13'h1210: data_buf = 8'h1f;
			13'h1211: data_buf = 8'h81;
			13'h1212: data_buf = 8'heb;
			13'h1213: data_buf = 8'hcd;
			13'h1214: data_buf = 8'hbd;
			13'h1215: data_buf = 8'h06;
			13'h1216: data_buf = 8'hca;
			13'h1217: data_buf = 8'h64;
			13'h1218: data_buf = 8'h12;
			13'h1219: data_buf = 8'hcd;
			13'h121a: data_buf = 8'heb;
			13'h121b: data_buf = 8'h16;
			13'h121c: data_buf = 8'h7b;
			13'h121d: data_buf = 8'he5;
			13'h121e: data_buf = 8'h09;
			13'h121f: data_buf = 8'hb7;
			13'h1220: data_buf = 8'hf2;
			13'h1221: data_buf = 8'h0d;
			13'h1222: data_buf = 8'h12;
			13'h1223: data_buf = 8'h22;
			13'h1224: data_buf = 8'h0a;
			13'h1225: data_buf = 8'h81;
			13'h1226: data_buf = 8'he1;
			13'h1227: data_buf = 8'h4e;
			13'h1228: data_buf = 8'h06;
			13'h1229: data_buf = 8'h00;
			13'h122a: data_buf = 8'h09;
			13'h122b: data_buf = 8'h09;
			13'h122c: data_buf = 8'h23;
			13'h122d: data_buf = 8'heb;
			13'h122e: data_buf = 8'h2a;
			13'h122f: data_buf = 8'h0a;
			13'h1230: data_buf = 8'h81;
			13'h1231: data_buf = 8'heb;
			13'h1232: data_buf = 8'hcd;
			13'h1233: data_buf = 8'hbd;
			13'h1234: data_buf = 8'h06;
			13'h1235: data_buf = 8'hca;
			13'h1236: data_buf = 8'h0e;
			13'h1237: data_buf = 8'h12;
			13'h1238: data_buf = 8'h01;
			13'h1239: data_buf = 8'h2d;
			13'h123a: data_buf = 8'h12;
			13'h123b: data_buf = 8'hc5;
			13'h123c: data_buf = 8'hf6;
			13'h123d: data_buf = 8'h80;
			13'h123e: data_buf = 8'h7e;
			13'h123f: data_buf = 8'h23;
			13'h1240: data_buf = 8'h23;
			13'h1241: data_buf = 8'h5e;
			13'h1242: data_buf = 8'h23;
			13'h1243: data_buf = 8'h56;
			13'h1244: data_buf = 8'h23;
			13'h1245: data_buf = 8'hf0;
			13'h1246: data_buf = 8'hb7;
			13'h1247: data_buf = 8'hc8;
			13'h1248: data_buf = 8'h44;
			13'h1249: data_buf = 8'h4d;
			13'h124a: data_buf = 8'h2a;
			13'h124b: data_buf = 8'h08;
			13'h124c: data_buf = 8'h81;
			13'h124d: data_buf = 8'hcd;
			13'h124e: data_buf = 8'hbd;
			13'h124f: data_buf = 8'h06;
			13'h1250: data_buf = 8'h60;
			13'h1251: data_buf = 8'h69;
			13'h1252: data_buf = 8'hd8;
			13'h1253: data_buf = 8'he1;
			13'h1254: data_buf = 8'he3;
			13'h1255: data_buf = 8'hcd;
			13'h1256: data_buf = 8'hbd;
			13'h1257: data_buf = 8'h06;
			13'h1258: data_buf = 8'he3;
			13'h1259: data_buf = 8'he5;
			13'h125a: data_buf = 8'h60;
			13'h125b: data_buf = 8'h69;
			13'h125c: data_buf = 8'hd0;
			13'h125d: data_buf = 8'hc1;
			13'h125e: data_buf = 8'hf1;
			13'h125f: data_buf = 8'hf1;
			13'h1260: data_buf = 8'he5;
			13'h1261: data_buf = 8'hd5;
			13'h1262: data_buf = 8'hc5;
			13'h1263: data_buf = 8'hc9;
			13'h1264: data_buf = 8'hd1;
			13'h1265: data_buf = 8'he1;
			13'h1266: data_buf = 8'h7d;
			13'h1267: data_buf = 8'hb4;
			13'h1268: data_buf = 8'hc8;
			13'h1269: data_buf = 8'h2b;
			13'h126a: data_buf = 8'h46;
			13'h126b: data_buf = 8'h2b;
			13'h126c: data_buf = 8'h4e;
			13'h126d: data_buf = 8'he5;
			13'h126e: data_buf = 8'h2b;
			13'h126f: data_buf = 8'h2b;
			13'h1270: data_buf = 8'h6e;
			13'h1271: data_buf = 8'h26;
			13'h1272: data_buf = 8'h00;
			13'h1273: data_buf = 8'h09;
			13'h1274: data_buf = 8'h50;
			13'h1275: data_buf = 8'h59;
			13'h1276: data_buf = 8'h2b;
			13'h1277: data_buf = 8'h44;
			13'h1278: data_buf = 8'h4d;
			13'h1279: data_buf = 8'h2a;
			13'h127a: data_buf = 8'h08;
			13'h127b: data_buf = 8'h81;
			13'h127c: data_buf = 8'hcd;
			13'h127d: data_buf = 8'hc4;
			13'h127e: data_buf = 8'h03;
			13'h127f: data_buf = 8'he1;
			13'h1280: data_buf = 8'h71;
			13'h1281: data_buf = 8'h23;
			13'h1282: data_buf = 8'h70;
			13'h1283: data_buf = 8'h69;
			13'h1284: data_buf = 8'h60;
			13'h1285: data_buf = 8'h2b;
			13'h1286: data_buf = 8'hc3;
			13'h1287: data_buf = 8'hd9;
			13'h1288: data_buf = 8'h11;
			13'h1289: data_buf = 8'hc5;
			13'h128a: data_buf = 8'he5;
			13'h128b: data_buf = 8'h2a;
			13'h128c: data_buf = 8'h29;
			13'h128d: data_buf = 8'h81;
			13'h128e: data_buf = 8'he3;
			13'h128f: data_buf = 8'hcd;
			13'h1290: data_buf = 8'h43;
			13'h1291: data_buf = 8'h0d;
			13'h1292: data_buf = 8'he3;
			13'h1293: data_buf = 8'hcd;
			13'h1294: data_buf = 8'hbe;
			13'h1295: data_buf = 8'h0c;
			13'h1296: data_buf = 8'h7e;
			13'h1297: data_buf = 8'he5;
			13'h1298: data_buf = 8'h2a;
			13'h1299: data_buf = 8'h29;
			13'h129a: data_buf = 8'h81;
			13'h129b: data_buf = 8'he5;
			13'h129c: data_buf = 8'h86;
			13'h129d: data_buf = 8'h1e;
			13'h129e: data_buf = 8'h1c;
			13'h129f: data_buf = 8'hda;
			13'h12a0: data_buf = 8'h09;
			13'h12a1: data_buf = 8'h04;
			13'h12a2: data_buf = 8'hcd;
			13'h12a3: data_buf = 8'h42;
			13'h12a4: data_buf = 8'h11;
			13'h12a5: data_buf = 8'hd1;
			13'h12a6: data_buf = 8'hcd;
			13'h12a7: data_buf = 8'hda;
			13'h12a8: data_buf = 8'h12;
			13'h12a9: data_buf = 8'he3;
			13'h12aa: data_buf = 8'hcd;
			13'h12ab: data_buf = 8'hd9;
			13'h12ac: data_buf = 8'h12;
			13'h12ad: data_buf = 8'he5;
			13'h12ae: data_buf = 8'h2a;
			13'h12af: data_buf = 8'h06;
			13'h12b0: data_buf = 8'h81;
			13'h12b1: data_buf = 8'heb;
			13'h12b2: data_buf = 8'hcd;
			13'h12b3: data_buf = 8'hc0;
			13'h12b4: data_buf = 8'h12;
			13'h12b5: data_buf = 8'hcd;
			13'h12b6: data_buf = 8'hc0;
			13'h12b7: data_buf = 8'h12;
			13'h12b8: data_buf = 8'h21;
			13'h12b9: data_buf = 8'hd8;
			13'h12ba: data_buf = 8'h0c;
			13'h12bb: data_buf = 8'he3;
			13'h12bc: data_buf = 8'he5;
			13'h12bd: data_buf = 8'hc3;
			13'h12be: data_buf = 8'h73;
			13'h12bf: data_buf = 8'h11;
			13'h12c0: data_buf = 8'he1;
			13'h12c1: data_buf = 8'he3;
			13'h12c2: data_buf = 8'h7e;
			13'h12c3: data_buf = 8'h23;
			13'h12c4: data_buf = 8'h23;
			13'h12c5: data_buf = 8'h4e;
			13'h12c6: data_buf = 8'h23;
			13'h12c7: data_buf = 8'h46;
			13'h12c8: data_buf = 8'h6f;
			13'h12c9: data_buf = 8'h2c;
			13'h12ca: data_buf = 8'h2d;
			13'h12cb: data_buf = 8'hc8;
			13'h12cc: data_buf = 8'h0a;
			13'h12cd: data_buf = 8'h12;
			13'h12ce: data_buf = 8'h03;
			13'h12cf: data_buf = 8'h13;
			13'h12d0: data_buf = 8'hc3;
			13'h12d1: data_buf = 8'hca;
			13'h12d2: data_buf = 8'h12;
			13'h12d3: data_buf = 8'hcd;
			13'h12d4: data_buf = 8'hbe;
			13'h12d5: data_buf = 8'h0c;
			13'h12d6: data_buf = 8'h2a;
			13'h12d7: data_buf = 8'h29;
			13'h12d8: data_buf = 8'h81;
			13'h12d9: data_buf = 8'heb;
			13'h12da: data_buf = 8'hcd;
			13'h12db: data_buf = 8'hf4;
			13'h12dc: data_buf = 8'h12;
			13'h12dd: data_buf = 8'heb;
			13'h12de: data_buf = 8'hc0;
			13'h12df: data_buf = 8'hd5;
			13'h12e0: data_buf = 8'h50;
			13'h12e1: data_buf = 8'h59;
			13'h12e2: data_buf = 8'h1b;
			13'h12e3: data_buf = 8'h4e;
			13'h12e4: data_buf = 8'h2a;
			13'h12e5: data_buf = 8'h08;
			13'h12e6: data_buf = 8'h81;
			13'h12e7: data_buf = 8'hcd;
			13'h12e8: data_buf = 8'hbd;
			13'h12e9: data_buf = 8'h06;
			13'h12ea: data_buf = 8'hc2;
			13'h12eb: data_buf = 8'hf2;
			13'h12ec: data_buf = 8'h12;
			13'h12ed: data_buf = 8'h47;
			13'h12ee: data_buf = 8'h09;
			13'h12ef: data_buf = 8'h22;
			13'h12f0: data_buf = 8'h08;
			13'h12f1: data_buf = 8'h81;
			13'h12f2: data_buf = 8'he1;
			13'h12f3: data_buf = 8'hc9;
			13'h12f4: data_buf = 8'h2a;
			13'h12f5: data_buf = 8'hf6;
			13'h12f6: data_buf = 8'h80;
			13'h12f7: data_buf = 8'h2b;
			13'h12f8: data_buf = 8'h46;
			13'h12f9: data_buf = 8'h2b;
			13'h12fa: data_buf = 8'h4e;
			13'h12fb: data_buf = 8'h2b;
			13'h12fc: data_buf = 8'h2b;
			13'h12fd: data_buf = 8'hcd;
			13'h12fe: data_buf = 8'hbd;
			13'h12ff: data_buf = 8'h06;
			13'h1300: data_buf = 8'hc0;
			13'h1301: data_buf = 8'h22;
			13'h1302: data_buf = 8'hf6;
			13'h1303: data_buf = 8'h80;
			13'h1304: data_buf = 8'hc9;
			13'h1305: data_buf = 8'h01;
			13'h1306: data_buf = 8'h84;
			13'h1307: data_buf = 8'h10;
			13'h1308: data_buf = 8'hc5;
			13'h1309: data_buf = 8'hcd;
			13'h130a: data_buf = 8'hd3;
			13'h130b: data_buf = 8'h12;
			13'h130c: data_buf = 8'haf;
			13'h130d: data_buf = 8'h57;
			13'h130e: data_buf = 8'h32;
			13'h130f: data_buf = 8'hf2;
			13'h1310: data_buf = 8'h80;
			13'h1311: data_buf = 8'h7e;
			13'h1312: data_buf = 8'hb7;
			13'h1313: data_buf = 8'hc9;
			13'h1314: data_buf = 8'h01;
			13'h1315: data_buf = 8'h84;
			13'h1316: data_buf = 8'h10;
			13'h1317: data_buf = 8'hc5;
			13'h1318: data_buf = 8'hcd;
			13'h1319: data_buf = 8'h09;
			13'h131a: data_buf = 8'h13;
			13'h131b: data_buf = 8'hca;
			13'h131c: data_buf = 8'h14;
			13'h131d: data_buf = 8'h09;
			13'h131e: data_buf = 8'h23;
			13'h131f: data_buf = 8'h23;
			13'h1320: data_buf = 8'h5e;
			13'h1321: data_buf = 8'h23;
			13'h1322: data_buf = 8'h56;
			13'h1323: data_buf = 8'h1a;
			13'h1324: data_buf = 8'hc9;
			13'h1325: data_buf = 8'h3e;
			13'h1326: data_buf = 8'h01;
			13'h1327: data_buf = 8'hcd;
			13'h1328: data_buf = 8'h42;
			13'h1329: data_buf = 8'h11;
			13'h132a: data_buf = 8'hcd;
			13'h132b: data_buf = 8'h1e;
			13'h132c: data_buf = 8'h14;
			13'h132d: data_buf = 8'h2a;
			13'h132e: data_buf = 8'h06;
			13'h132f: data_buf = 8'h81;
			13'h1330: data_buf = 8'h73;
			13'h1331: data_buf = 8'hc1;
			13'h1332: data_buf = 8'hc3;
			13'h1333: data_buf = 8'h73;
			13'h1334: data_buf = 8'h11;
			13'h1335: data_buf = 8'hcd;
			13'h1336: data_buf = 8'hce;
			13'h1337: data_buf = 8'h13;
			13'h1338: data_buf = 8'haf;
			13'h1339: data_buf = 8'he3;
			13'h133a: data_buf = 8'h4f;
			13'h133b: data_buf = 8'he5;
			13'h133c: data_buf = 8'h7e;
			13'h133d: data_buf = 8'hb8;
			13'h133e: data_buf = 8'hda;
			13'h133f: data_buf = 8'h43;
			13'h1340: data_buf = 8'h13;
			13'h1341: data_buf = 8'h78;
			13'h1342: data_buf = 8'h11;
			13'h1343: data_buf = 8'h0e;
			13'h1344: data_buf = 8'h00;
			13'h1345: data_buf = 8'hc5;
			13'h1346: data_buf = 8'hcd;
			13'h1347: data_buf = 8'hac;
			13'h1348: data_buf = 8'h11;
			13'h1349: data_buf = 8'hc1;
			13'h134a: data_buf = 8'he1;
			13'h134b: data_buf = 8'he5;
			13'h134c: data_buf = 8'h23;
			13'h134d: data_buf = 8'h23;
			13'h134e: data_buf = 8'h46;
			13'h134f: data_buf = 8'h23;
			13'h1350: data_buf = 8'h66;
			13'h1351: data_buf = 8'h68;
			13'h1352: data_buf = 8'h06;
			13'h1353: data_buf = 8'h00;
			13'h1354: data_buf = 8'h09;
			13'h1355: data_buf = 8'h44;
			13'h1356: data_buf = 8'h4d;
			13'h1357: data_buf = 8'hcd;
			13'h1358: data_buf = 8'h45;
			13'h1359: data_buf = 8'h11;
			13'h135a: data_buf = 8'h6f;
			13'h135b: data_buf = 8'hcd;
			13'h135c: data_buf = 8'hc9;
			13'h135d: data_buf = 8'h12;
			13'h135e: data_buf = 8'hd1;
			13'h135f: data_buf = 8'hcd;
			13'h1360: data_buf = 8'hda;
			13'h1361: data_buf = 8'h12;
			13'h1362: data_buf = 8'hc3;
			13'h1363: data_buf = 8'h73;
			13'h1364: data_buf = 8'h11;
			13'h1365: data_buf = 8'hcd;
			13'h1366: data_buf = 8'hce;
			13'h1367: data_buf = 8'h13;
			13'h1368: data_buf = 8'hd1;
			13'h1369: data_buf = 8'hd5;
			13'h136a: data_buf = 8'h1a;
			13'h136b: data_buf = 8'h90;
			13'h136c: data_buf = 8'hc3;
			13'h136d: data_buf = 8'h39;
			13'h136e: data_buf = 8'h13;
			13'h136f: data_buf = 8'heb;
			13'h1370: data_buf = 8'h7e;
			13'h1371: data_buf = 8'hcd;
			13'h1372: data_buf = 8'hd3;
			13'h1373: data_buf = 8'h13;
			13'h1374: data_buf = 8'h04;
			13'h1375: data_buf = 8'h05;
			13'h1376: data_buf = 8'hca;
			13'h1377: data_buf = 8'h14;
			13'h1378: data_buf = 8'h09;
			13'h1379: data_buf = 8'hc5;
			13'h137a: data_buf = 8'h1e;
			13'h137b: data_buf = 8'hff;
			13'h137c: data_buf = 8'hfe;
			13'h137d: data_buf = 8'h29;
			13'h137e: data_buf = 8'hca;
			13'h137f: data_buf = 8'h88;
			13'h1380: data_buf = 8'h13;
			13'h1381: data_buf = 8'hcd;
			13'h1382: data_buf = 8'hc3;
			13'h1383: data_buf = 8'h06;
			13'h1384: data_buf = 8'h2c;
			13'h1385: data_buf = 8'hcd;
			13'h1386: data_buf = 8'h1b;
			13'h1387: data_buf = 8'h14;
			13'h1388: data_buf = 8'hcd;
			13'h1389: data_buf = 8'hc3;
			13'h138a: data_buf = 8'h06;
			13'h138b: data_buf = 8'h29;
			13'h138c: data_buf = 8'hf1;
			13'h138d: data_buf = 8'he3;
			13'h138e: data_buf = 8'h01;
			13'h138f: data_buf = 8'h3b;
			13'h1390: data_buf = 8'h13;
			13'h1391: data_buf = 8'hc5;
			13'h1392: data_buf = 8'h3d;
			13'h1393: data_buf = 8'hbe;
			13'h1394: data_buf = 8'h06;
			13'h1395: data_buf = 8'h00;
			13'h1396: data_buf = 8'hd0;
			13'h1397: data_buf = 8'h4f;
			13'h1398: data_buf = 8'h7e;
			13'h1399: data_buf = 8'h91;
			13'h139a: data_buf = 8'hbb;
			13'h139b: data_buf = 8'h47;
			13'h139c: data_buf = 8'hd8;
			13'h139d: data_buf = 8'h43;
			13'h139e: data_buf = 8'hc9;
			13'h139f: data_buf = 8'hcd;
			13'h13a0: data_buf = 8'h09;
			13'h13a1: data_buf = 8'h13;
			13'h13a2: data_buf = 8'hca;
			13'h13a3: data_buf = 8'hbc;
			13'h13a4: data_buf = 8'h14;
			13'h13a5: data_buf = 8'h5f;
			13'h13a6: data_buf = 8'h23;
			13'h13a7: data_buf = 8'h23;
			13'h13a8: data_buf = 8'h7e;
			13'h13a9: data_buf = 8'h23;
			13'h13aa: data_buf = 8'h66;
			13'h13ab: data_buf = 8'h6f;
			13'h13ac: data_buf = 8'he5;
			13'h13ad: data_buf = 8'h19;
			13'h13ae: data_buf = 8'h46;
			13'h13af: data_buf = 8'h72;
			13'h13b0: data_buf = 8'he3;
			13'h13b1: data_buf = 8'hc5;
			13'h13b2: data_buf = 8'h7e;
			13'h13b3: data_buf = 8'hfe;
			13'h13b4: data_buf = 8'h24;
			13'h13b5: data_buf = 8'hc2;
			13'h13b6: data_buf = 8'hbd;
			13'h13b7: data_buf = 8'h13;
			13'h13b8: data_buf = 8'hcd;
			13'h13b9: data_buf = 8'he7;
			13'h13ba: data_buf = 8'h1b;
			13'h13bb: data_buf = 8'h18;
			13'h13bc: data_buf = 8'h0d;
			13'h13bd: data_buf = 8'hfe;
			13'h13be: data_buf = 8'h25;
			13'h13bf: data_buf = 8'hc2;
			13'h13c0: data_buf = 8'hc7;
			13'h13c1: data_buf = 8'h13;
			13'h13c2: data_buf = 8'hcd;
			13'h13c3: data_buf = 8'h57;
			13'h13c4: data_buf = 8'h1c;
			13'h13c5: data_buf = 8'h18;
			13'h13c6: data_buf = 8'h03;
			13'h13c7: data_buf = 8'hcd;
			13'h13c8: data_buf = 8'ha3;
			13'h13c9: data_buf = 8'h17;
			13'h13ca: data_buf = 8'hc1;
			13'h13cb: data_buf = 8'he1;
			13'h13cc: data_buf = 8'h70;
			13'h13cd: data_buf = 8'hc9;
			13'h13ce: data_buf = 8'heb;
			13'h13cf: data_buf = 8'hcd;
			13'h13d0: data_buf = 8'hc3;
			13'h13d1: data_buf = 8'h06;
			13'h13d2: data_buf = 8'h29;
			13'h13d3: data_buf = 8'hc1;
			13'h13d4: data_buf = 8'hd1;
			13'h13d5: data_buf = 8'hc5;
			13'h13d6: data_buf = 8'h43;
			13'h13d7: data_buf = 8'hc9;
			13'h13d8: data_buf = 8'hcd;
			13'h13d9: data_buf = 8'h1e;
			13'h13da: data_buf = 8'h14;
			13'h13db: data_buf = 8'h32;
			13'h13dc: data_buf = 8'h84;
			13'h13dd: data_buf = 8'h80;
			13'h13de: data_buf = 8'hcd;
			13'h13df: data_buf = 8'h83;
			13'h13e0: data_buf = 8'h80;
			13'h13e1: data_buf = 8'hc3;
			13'h13e2: data_buf = 8'h84;
			13'h13e3: data_buf = 8'h10;
			13'h13e4: data_buf = 8'hcd;
			13'h13e5: data_buf = 8'h08;
			13'h13e6: data_buf = 8'h14;
			13'h13e7: data_buf = 8'hc3;
			13'h13e8: data_buf = 8'h4b;
			13'h13e9: data_buf = 8'h80;
			13'h13ea: data_buf = 8'hcd;
			13'h13eb: data_buf = 8'h08;
			13'h13ec: data_buf = 8'h14;
			13'h13ed: data_buf = 8'hf5;
			13'h13ee: data_buf = 8'h1e;
			13'h13ef: data_buf = 8'h00;
			13'h13f0: data_buf = 8'h2b;
			13'h13f1: data_buf = 8'hcd;
			13'h13f2: data_buf = 8'h4d;
			13'h13f3: data_buf = 8'h08;
			13'h13f4: data_buf = 8'hca;
			13'h13f5: data_buf = 8'hfe;
			13'h13f6: data_buf = 8'h13;
			13'h13f7: data_buf = 8'hcd;
			13'h13f8: data_buf = 8'hc3;
			13'h13f9: data_buf = 8'h06;
			13'h13fa: data_buf = 8'h2c;
			13'h13fb: data_buf = 8'hcd;
			13'h13fc: data_buf = 8'h1b;
			13'h13fd: data_buf = 8'h14;
			13'h13fe: data_buf = 8'hc1;
			13'h13ff: data_buf = 8'hcd;
			13'h1400: data_buf = 8'h83;
			13'h1401: data_buf = 8'h80;
			13'h1402: data_buf = 8'hab;
			13'h1403: data_buf = 8'ha0;
			13'h1404: data_buf = 8'hca;
			13'h1405: data_buf = 8'hff;
			13'h1406: data_buf = 8'h13;
			13'h1407: data_buf = 8'hc9;
			13'h1408: data_buf = 8'hcd;
			13'h1409: data_buf = 8'h1b;
			13'h140a: data_buf = 8'h14;
			13'h140b: data_buf = 8'h32;
			13'h140c: data_buf = 8'h84;
			13'h140d: data_buf = 8'h80;
			13'h140e: data_buf = 8'h32;
			13'h140f: data_buf = 8'h4c;
			13'h1410: data_buf = 8'h80;
			13'h1411: data_buf = 8'hcd;
			13'h1412: data_buf = 8'hc3;
			13'h1413: data_buf = 8'h06;
			13'h1414: data_buf = 8'h2c;
			13'h1415: data_buf = 8'hc3;
			13'h1416: data_buf = 8'h1b;
			13'h1417: data_buf = 8'h14;
			13'h1418: data_buf = 8'hcd;
			13'h1419: data_buf = 8'h4d;
			13'h141a: data_buf = 8'h08;
			13'h141b: data_buf = 8'hcd;
			13'h141c: data_buf = 8'hba;
			13'h141d: data_buf = 8'h0c;
			13'h141e: data_buf = 8'hcd;
			13'h141f: data_buf = 8'hf9;
			13'h1420: data_buf = 8'h08;
			13'h1421: data_buf = 8'h7a;
			13'h1422: data_buf = 8'hb7;
			13'h1423: data_buf = 8'hc2;
			13'h1424: data_buf = 8'h14;
			13'h1425: data_buf = 8'h09;
			13'h1426: data_buf = 8'h2b;
			13'h1427: data_buf = 8'hcd;
			13'h1428: data_buf = 8'h4d;
			13'h1429: data_buf = 8'h08;
			13'h142a: data_buf = 8'h7b;
			13'h142b: data_buf = 8'hc9;
			13'h142c: data_buf = 8'hcd;
			13'h142d: data_buf = 8'hff;
			13'h142e: data_buf = 8'h08;
			13'h142f: data_buf = 8'h1a;
			13'h1430: data_buf = 8'hc3;
			13'h1431: data_buf = 8'h84;
			13'h1432: data_buf = 8'h10;
			13'h1433: data_buf = 8'hcd;
			13'h1434: data_buf = 8'hba;
			13'h1435: data_buf = 8'h0c;
			13'h1436: data_buf = 8'hcd;
			13'h1437: data_buf = 8'hff;
			13'h1438: data_buf = 8'h08;
			13'h1439: data_buf = 8'hd5;
			13'h143a: data_buf = 8'hcd;
			13'h143b: data_buf = 8'hc3;
			13'h143c: data_buf = 8'h06;
			13'h143d: data_buf = 8'h2c;
			13'h143e: data_buf = 8'hcd;
			13'h143f: data_buf = 8'h1b;
			13'h1440: data_buf = 8'h14;
			13'h1441: data_buf = 8'hd1;
			13'h1442: data_buf = 8'h12;
			13'h1443: data_buf = 8'hc9;
			13'h1444: data_buf = 8'h21;
			13'h1445: data_buf = 8'h1a;
			13'h1446: data_buf = 8'h19;
			13'h1447: data_buf = 8'hcd;
			13'h1448: data_buf = 8'heb;
			13'h1449: data_buf = 8'h16;
			13'h144a: data_buf = 8'hc3;
			13'h144b: data_buf = 8'h56;
			13'h144c: data_buf = 8'h14;
			13'h144d: data_buf = 8'hcd;
			13'h144e: data_buf = 8'heb;
			13'h144f: data_buf = 8'h16;
			13'h1450: data_buf = 8'h21;
			13'h1451: data_buf = 8'hc1;
			13'h1452: data_buf = 8'hd1;
			13'h1453: data_buf = 8'hcd;
			13'h1454: data_buf = 8'hc5;
			13'h1455: data_buf = 8'h16;
			13'h1456: data_buf = 8'h78;
			13'h1457: data_buf = 8'hb7;
			13'h1458: data_buf = 8'hc8;
			13'h1459: data_buf = 8'h3a;
			13'h145a: data_buf = 8'h2c;
			13'h145b: data_buf = 8'h81;
			13'h145c: data_buf = 8'hb7;
			13'h145d: data_buf = 8'hca;
			13'h145e: data_buf = 8'hdd;
			13'h145f: data_buf = 8'h16;
			13'h1460: data_buf = 8'h90;
			13'h1461: data_buf = 8'hd2;
			13'h1462: data_buf = 8'h70;
			13'h1463: data_buf = 8'h14;
			13'h1464: data_buf = 8'h2f;
			13'h1465: data_buf = 8'h3c;
			13'h1466: data_buf = 8'heb;
			13'h1467: data_buf = 8'hcd;
			13'h1468: data_buf = 8'hcd;
			13'h1469: data_buf = 8'h16;
			13'h146a: data_buf = 8'heb;
			13'h146b: data_buf = 8'hcd;
			13'h146c: data_buf = 8'hdd;
			13'h146d: data_buf = 8'h16;
			13'h146e: data_buf = 8'hc1;
			13'h146f: data_buf = 8'hd1;
			13'h1470: data_buf = 8'hfe;
			13'h1471: data_buf = 8'h19;
			13'h1472: data_buf = 8'hd0;
			13'h1473: data_buf = 8'hf5;
			13'h1474: data_buf = 8'hcd;
			13'h1475: data_buf = 8'h02;
			13'h1476: data_buf = 8'h17;
			13'h1477: data_buf = 8'h67;
			13'h1478: data_buf = 8'hf1;
			13'h1479: data_buf = 8'hcd;
			13'h147a: data_buf = 8'h1b;
			13'h147b: data_buf = 8'h15;
			13'h147c: data_buf = 8'hb4;
			13'h147d: data_buf = 8'h21;
			13'h147e: data_buf = 8'h29;
			13'h147f: data_buf = 8'h81;
			13'h1480: data_buf = 8'hf2;
			13'h1481: data_buf = 8'h96;
			13'h1482: data_buf = 8'h14;
			13'h1483: data_buf = 8'hcd;
			13'h1484: data_buf = 8'hfb;
			13'h1485: data_buf = 8'h14;
			13'h1486: data_buf = 8'hd2;
			13'h1487: data_buf = 8'hdc;
			13'h1488: data_buf = 8'h14;
			13'h1489: data_buf = 8'h23;
			13'h148a: data_buf = 8'h34;
			13'h148b: data_buf = 8'hca;
			13'h148c: data_buf = 8'h04;
			13'h148d: data_buf = 8'h04;
			13'h148e: data_buf = 8'h2e;
			13'h148f: data_buf = 8'h01;
			13'h1490: data_buf = 8'hcd;
			13'h1491: data_buf = 8'h31;
			13'h1492: data_buf = 8'h15;
			13'h1493: data_buf = 8'hc3;
			13'h1494: data_buf = 8'hdc;
			13'h1495: data_buf = 8'h14;
			13'h1496: data_buf = 8'haf;
			13'h1497: data_buf = 8'h90;
			13'h1498: data_buf = 8'h47;
			13'h1499: data_buf = 8'h7e;
			13'h149a: data_buf = 8'h9b;
			13'h149b: data_buf = 8'h5f;
			13'h149c: data_buf = 8'h23;
			13'h149d: data_buf = 8'h7e;
			13'h149e: data_buf = 8'h9a;
			13'h149f: data_buf = 8'h57;
			13'h14a0: data_buf = 8'h23;
			13'h14a1: data_buf = 8'h7e;
			13'h14a2: data_buf = 8'h99;
			13'h14a3: data_buf = 8'h4f;
			13'h14a4: data_buf = 8'hdc;
			13'h14a5: data_buf = 8'h07;
			13'h14a6: data_buf = 8'h15;
			13'h14a7: data_buf = 8'h68;
			13'h14a8: data_buf = 8'h63;
			13'h14a9: data_buf = 8'haf;
			13'h14aa: data_buf = 8'h47;
			13'h14ab: data_buf = 8'h79;
			13'h14ac: data_buf = 8'hb7;
			13'h14ad: data_buf = 8'hc2;
			13'h14ae: data_buf = 8'hc9;
			13'h14af: data_buf = 8'h14;
			13'h14b0: data_buf = 8'h4a;
			13'h14b1: data_buf = 8'h54;
			13'h14b2: data_buf = 8'h65;
			13'h14b3: data_buf = 8'h6f;
			13'h14b4: data_buf = 8'h78;
			13'h14b5: data_buf = 8'hd6;
			13'h14b6: data_buf = 8'h08;
			13'h14b7: data_buf = 8'hfe;
			13'h14b8: data_buf = 8'he0;
			13'h14b9: data_buf = 8'hc2;
			13'h14ba: data_buf = 8'haa;
			13'h14bb: data_buf = 8'h14;
			13'h14bc: data_buf = 8'haf;
			13'h14bd: data_buf = 8'h32;
			13'h14be: data_buf = 8'h2c;
			13'h14bf: data_buf = 8'h81;
			13'h14c0: data_buf = 8'hc9;
			13'h14c1: data_buf = 8'h05;
			13'h14c2: data_buf = 8'h29;
			13'h14c3: data_buf = 8'h7a;
			13'h14c4: data_buf = 8'h17;
			13'h14c5: data_buf = 8'h57;
			13'h14c6: data_buf = 8'h79;
			13'h14c7: data_buf = 8'h8f;
			13'h14c8: data_buf = 8'h4f;
			13'h14c9: data_buf = 8'hf2;
			13'h14ca: data_buf = 8'hc1;
			13'h14cb: data_buf = 8'h14;
			13'h14cc: data_buf = 8'h78;
			13'h14cd: data_buf = 8'h5c;
			13'h14ce: data_buf = 8'h45;
			13'h14cf: data_buf = 8'hb7;
			13'h14d0: data_buf = 8'hca;
			13'h14d1: data_buf = 8'hdc;
			13'h14d2: data_buf = 8'h14;
			13'h14d3: data_buf = 8'h21;
			13'h14d4: data_buf = 8'h2c;
			13'h14d5: data_buf = 8'h81;
			13'h14d6: data_buf = 8'h86;
			13'h14d7: data_buf = 8'h77;
			13'h14d8: data_buf = 8'hd2;
			13'h14d9: data_buf = 8'hbc;
			13'h14da: data_buf = 8'h14;
			13'h14db: data_buf = 8'hc8;
			13'h14dc: data_buf = 8'h78;
			13'h14dd: data_buf = 8'h21;
			13'h14de: data_buf = 8'h2c;
			13'h14df: data_buf = 8'h81;
			13'h14e0: data_buf = 8'hb7;
			13'h14e1: data_buf = 8'hfc;
			13'h14e2: data_buf = 8'hee;
			13'h14e3: data_buf = 8'h14;
			13'h14e4: data_buf = 8'h46;
			13'h14e5: data_buf = 8'h23;
			13'h14e6: data_buf = 8'h7e;
			13'h14e7: data_buf = 8'he6;
			13'h14e8: data_buf = 8'h80;
			13'h14e9: data_buf = 8'ha9;
			13'h14ea: data_buf = 8'h4f;
			13'h14eb: data_buf = 8'hc3;
			13'h14ec: data_buf = 8'hdd;
			13'h14ed: data_buf = 8'h16;
			13'h14ee: data_buf = 8'h1c;
			13'h14ef: data_buf = 8'hc0;
			13'h14f0: data_buf = 8'h14;
			13'h14f1: data_buf = 8'hc0;
			13'h14f2: data_buf = 8'h0c;
			13'h14f3: data_buf = 8'hc0;
			13'h14f4: data_buf = 8'h0e;
			13'h14f5: data_buf = 8'h80;
			13'h14f6: data_buf = 8'h34;
			13'h14f7: data_buf = 8'hc0;
			13'h14f8: data_buf = 8'hc3;
			13'h14f9: data_buf = 8'h04;
			13'h14fa: data_buf = 8'h04;
			13'h14fb: data_buf = 8'h7e;
			13'h14fc: data_buf = 8'h83;
			13'h14fd: data_buf = 8'h5f;
			13'h14fe: data_buf = 8'h23;
			13'h14ff: data_buf = 8'h7e;
			13'h1500: data_buf = 8'h8a;
			13'h1501: data_buf = 8'h57;
			13'h1502: data_buf = 8'h23;
			13'h1503: data_buf = 8'h7e;
			13'h1504: data_buf = 8'h89;
			13'h1505: data_buf = 8'h4f;
			13'h1506: data_buf = 8'hc9;
			13'h1507: data_buf = 8'h21;
			13'h1508: data_buf = 8'h2d;
			13'h1509: data_buf = 8'h81;
			13'h150a: data_buf = 8'h7e;
			13'h150b: data_buf = 8'h2f;
			13'h150c: data_buf = 8'h77;
			13'h150d: data_buf = 8'haf;
			13'h150e: data_buf = 8'h6f;
			13'h150f: data_buf = 8'h90;
			13'h1510: data_buf = 8'h47;
			13'h1511: data_buf = 8'h7d;
			13'h1512: data_buf = 8'h9b;
			13'h1513: data_buf = 8'h5f;
			13'h1514: data_buf = 8'h7d;
			13'h1515: data_buf = 8'h9a;
			13'h1516: data_buf = 8'h57;
			13'h1517: data_buf = 8'h7d;
			13'h1518: data_buf = 8'h99;
			13'h1519: data_buf = 8'h4f;
			13'h151a: data_buf = 8'hc9;
			13'h151b: data_buf = 8'h06;
			13'h151c: data_buf = 8'h00;
			13'h151d: data_buf = 8'hd6;
			13'h151e: data_buf = 8'h08;
			13'h151f: data_buf = 8'hda;
			13'h1520: data_buf = 8'h2a;
			13'h1521: data_buf = 8'h15;
			13'h1522: data_buf = 8'h43;
			13'h1523: data_buf = 8'h5a;
			13'h1524: data_buf = 8'h51;
			13'h1525: data_buf = 8'h0e;
			13'h1526: data_buf = 8'h00;
			13'h1527: data_buf = 8'hc3;
			13'h1528: data_buf = 8'h1d;
			13'h1529: data_buf = 8'h15;
			13'h152a: data_buf = 8'hc6;
			13'h152b: data_buf = 8'h09;
			13'h152c: data_buf = 8'h6f;
			13'h152d: data_buf = 8'haf;
			13'h152e: data_buf = 8'h2d;
			13'h152f: data_buf = 8'hc8;
			13'h1530: data_buf = 8'h79;
			13'h1531: data_buf = 8'h1f;
			13'h1532: data_buf = 8'h4f;
			13'h1533: data_buf = 8'h7a;
			13'h1534: data_buf = 8'h1f;
			13'h1535: data_buf = 8'h57;
			13'h1536: data_buf = 8'h7b;
			13'h1537: data_buf = 8'h1f;
			13'h1538: data_buf = 8'h5f;
			13'h1539: data_buf = 8'h78;
			13'h153a: data_buf = 8'h1f;
			13'h153b: data_buf = 8'h47;
			13'h153c: data_buf = 8'hc3;
			13'h153d: data_buf = 8'h2d;
			13'h153e: data_buf = 8'h15;
			13'h153f: data_buf = 8'h00;
			13'h1540: data_buf = 8'h00;
			13'h1541: data_buf = 8'h00;
			13'h1542: data_buf = 8'h81;
			13'h1543: data_buf = 8'h03;
			13'h1544: data_buf = 8'haa;
			13'h1545: data_buf = 8'h56;
			13'h1546: data_buf = 8'h19;
			13'h1547: data_buf = 8'h80;
			13'h1548: data_buf = 8'hf1;
			13'h1549: data_buf = 8'h22;
			13'h154a: data_buf = 8'h76;
			13'h154b: data_buf = 8'h80;
			13'h154c: data_buf = 8'h45;
			13'h154d: data_buf = 8'haa;
			13'h154e: data_buf = 8'h38;
			13'h154f: data_buf = 8'h82;
			13'h1550: data_buf = 8'hcd;
			13'h1551: data_buf = 8'h9c;
			13'h1552: data_buf = 8'h16;
			13'h1553: data_buf = 8'hb7;
			13'h1554: data_buf = 8'hea;
			13'h1555: data_buf = 8'h14;
			13'h1556: data_buf = 8'h09;
			13'h1557: data_buf = 8'h21;
			13'h1558: data_buf = 8'h2c;
			13'h1559: data_buf = 8'h81;
			13'h155a: data_buf = 8'h7e;
			13'h155b: data_buf = 8'h01;
			13'h155c: data_buf = 8'h35;
			13'h155d: data_buf = 8'h80;
			13'h155e: data_buf = 8'h11;
			13'h155f: data_buf = 8'hf3;
			13'h1560: data_buf = 8'h04;
			13'h1561: data_buf = 8'h90;
			13'h1562: data_buf = 8'hf5;
			13'h1563: data_buf = 8'h70;
			13'h1564: data_buf = 8'hd5;
			13'h1565: data_buf = 8'hc5;
			13'h1566: data_buf = 8'hcd;
			13'h1567: data_buf = 8'h56;
			13'h1568: data_buf = 8'h14;
			13'h1569: data_buf = 8'hc1;
			13'h156a: data_buf = 8'hd1;
			13'h156b: data_buf = 8'h04;
			13'h156c: data_buf = 8'hcd;
			13'h156d: data_buf = 8'hf2;
			13'h156e: data_buf = 8'h15;
			13'h156f: data_buf = 8'h21;
			13'h1570: data_buf = 8'h3f;
			13'h1571: data_buf = 8'h15;
			13'h1572: data_buf = 8'hcd;
			13'h1573: data_buf = 8'h4d;
			13'h1574: data_buf = 8'h14;
			13'h1575: data_buf = 8'h21;
			13'h1576: data_buf = 8'h43;
			13'h1577: data_buf = 8'h15;
			13'h1578: data_buf = 8'hcd;
			13'h1579: data_buf = 8'he4;
			13'h157a: data_buf = 8'h19;
			13'h157b: data_buf = 8'h01;
			13'h157c: data_buf = 8'h80;
			13'h157d: data_buf = 8'h80;
			13'h157e: data_buf = 8'h11;
			13'h157f: data_buf = 8'h00;
			13'h1580: data_buf = 8'h00;
			13'h1581: data_buf = 8'hcd;
			13'h1582: data_buf = 8'h56;
			13'h1583: data_buf = 8'h14;
			13'h1584: data_buf = 8'hf1;
			13'h1585: data_buf = 8'hcd;
			13'h1586: data_buf = 8'h17;
			13'h1587: data_buf = 8'h18;
			13'h1588: data_buf = 8'h01;
			13'h1589: data_buf = 8'h31;
			13'h158a: data_buf = 8'h80;
			13'h158b: data_buf = 8'h11;
			13'h158c: data_buf = 8'h18;
			13'h158d: data_buf = 8'h72;
			13'h158e: data_buf = 8'h21;
			13'h158f: data_buf = 8'hc1;
			13'h1590: data_buf = 8'hd1;
			13'h1591: data_buf = 8'hcd;
			13'h1592: data_buf = 8'h9c;
			13'h1593: data_buf = 8'h16;
			13'h1594: data_buf = 8'hc8;
			13'h1595: data_buf = 8'h2e;
			13'h1596: data_buf = 8'h00;
			13'h1597: data_buf = 8'hcd;
			13'h1598: data_buf = 8'h5a;
			13'h1599: data_buf = 8'h16;
			13'h159a: data_buf = 8'h79;
			13'h159b: data_buf = 8'h32;
			13'h159c: data_buf = 8'h3b;
			13'h159d: data_buf = 8'h81;
			13'h159e: data_buf = 8'heb;
			13'h159f: data_buf = 8'h22;
			13'h15a0: data_buf = 8'h3c;
			13'h15a1: data_buf = 8'h81;
			13'h15a2: data_buf = 8'h01;
			13'h15a3: data_buf = 8'h00;
			13'h15a4: data_buf = 8'h00;
			13'h15a5: data_buf = 8'h50;
			13'h15a6: data_buf = 8'h58;
			13'h15a7: data_buf = 8'h21;
			13'h15a8: data_buf = 8'ha7;
			13'h15a9: data_buf = 8'h14;
			13'h15aa: data_buf = 8'he5;
			13'h15ab: data_buf = 8'h21;
			13'h15ac: data_buf = 8'hb3;
			13'h15ad: data_buf = 8'h15;
			13'h15ae: data_buf = 8'he5;
			13'h15af: data_buf = 8'he5;
			13'h15b0: data_buf = 8'h21;
			13'h15b1: data_buf = 8'h29;
			13'h15b2: data_buf = 8'h81;
			13'h15b3: data_buf = 8'h7e;
			13'h15b4: data_buf = 8'h23;
			13'h15b5: data_buf = 8'hb7;
			13'h15b6: data_buf = 8'hca;
			13'h15b7: data_buf = 8'hdf;
			13'h15b8: data_buf = 8'h15;
			13'h15b9: data_buf = 8'he5;
			13'h15ba: data_buf = 8'h2e;
			13'h15bb: data_buf = 8'h08;
			13'h15bc: data_buf = 8'h1f;
			13'h15bd: data_buf = 8'h67;
			13'h15be: data_buf = 8'h79;
			13'h15bf: data_buf = 8'hd2;
			13'h15c0: data_buf = 8'hcd;
			13'h15c1: data_buf = 8'h15;
			13'h15c2: data_buf = 8'he5;
			13'h15c3: data_buf = 8'h2a;
			13'h15c4: data_buf = 8'h3c;
			13'h15c5: data_buf = 8'h81;
			13'h15c6: data_buf = 8'h19;
			13'h15c7: data_buf = 8'heb;
			13'h15c8: data_buf = 8'he1;
			13'h15c9: data_buf = 8'h3a;
			13'h15ca: data_buf = 8'h3b;
			13'h15cb: data_buf = 8'h81;
			13'h15cc: data_buf = 8'h89;
			13'h15cd: data_buf = 8'h1f;
			13'h15ce: data_buf = 8'h4f;
			13'h15cf: data_buf = 8'h7a;
			13'h15d0: data_buf = 8'h1f;
			13'h15d1: data_buf = 8'h57;
			13'h15d2: data_buf = 8'h7b;
			13'h15d3: data_buf = 8'h1f;
			13'h15d4: data_buf = 8'h5f;
			13'h15d5: data_buf = 8'h78;
			13'h15d6: data_buf = 8'h1f;
			13'h15d7: data_buf = 8'h47;
			13'h15d8: data_buf = 8'h2d;
			13'h15d9: data_buf = 8'h7c;
			13'h15da: data_buf = 8'hc2;
			13'h15db: data_buf = 8'hbc;
			13'h15dc: data_buf = 8'h15;
			13'h15dd: data_buf = 8'he1;
			13'h15de: data_buf = 8'hc9;
			13'h15df: data_buf = 8'h43;
			13'h15e0: data_buf = 8'h5a;
			13'h15e1: data_buf = 8'h51;
			13'h15e2: data_buf = 8'h4f;
			13'h15e3: data_buf = 8'hc9;
			13'h15e4: data_buf = 8'hcd;
			13'h15e5: data_buf = 8'hcd;
			13'h15e6: data_buf = 8'h16;
			13'h15e7: data_buf = 8'h01;
			13'h15e8: data_buf = 8'h20;
			13'h15e9: data_buf = 8'h84;
			13'h15ea: data_buf = 8'h11;
			13'h15eb: data_buf = 8'h00;
			13'h15ec: data_buf = 8'h00;
			13'h15ed: data_buf = 8'hcd;
			13'h15ee: data_buf = 8'hdd;
			13'h15ef: data_buf = 8'h16;
			13'h15f0: data_buf = 8'hc1;
			13'h15f1: data_buf = 8'hd1;
			13'h15f2: data_buf = 8'hcd;
			13'h15f3: data_buf = 8'h9c;
			13'h15f4: data_buf = 8'h16;
			13'h15f5: data_buf = 8'hca;
			13'h15f6: data_buf = 8'hf8;
			13'h15f7: data_buf = 8'h03;
			13'h15f8: data_buf = 8'h2e;
			13'h15f9: data_buf = 8'hff;
			13'h15fa: data_buf = 8'hcd;
			13'h15fb: data_buf = 8'h5a;
			13'h15fc: data_buf = 8'h16;
			13'h15fd: data_buf = 8'h34;
			13'h15fe: data_buf = 8'h34;
			13'h15ff: data_buf = 8'h2b;
			13'h1600: data_buf = 8'h7e;
			13'h1601: data_buf = 8'h32;
			13'h1602: data_buf = 8'h57;
			13'h1603: data_buf = 8'h80;
			13'h1604: data_buf = 8'h2b;
			13'h1605: data_buf = 8'h7e;
			13'h1606: data_buf = 8'h32;
			13'h1607: data_buf = 8'h53;
			13'h1608: data_buf = 8'h80;
			13'h1609: data_buf = 8'h2b;
			13'h160a: data_buf = 8'h7e;
			13'h160b: data_buf = 8'h32;
			13'h160c: data_buf = 8'h4f;
			13'h160d: data_buf = 8'h80;
			13'h160e: data_buf = 8'h41;
			13'h160f: data_buf = 8'heb;
			13'h1610: data_buf = 8'haf;
			13'h1611: data_buf = 8'h4f;
			13'h1612: data_buf = 8'h57;
			13'h1613: data_buf = 8'h5f;
			13'h1614: data_buf = 8'h32;
			13'h1615: data_buf = 8'h5a;
			13'h1616: data_buf = 8'h80;
			13'h1617: data_buf = 8'he5;
			13'h1618: data_buf = 8'hc5;
			13'h1619: data_buf = 8'h7d;
			13'h161a: data_buf = 8'hcd;
			13'h161b: data_buf = 8'h4e;
			13'h161c: data_buf = 8'h80;
			13'h161d: data_buf = 8'hde;
			13'h161e: data_buf = 8'h00;
			13'h161f: data_buf = 8'h3f;
			13'h1620: data_buf = 8'hd2;
			13'h1621: data_buf = 8'h2a;
			13'h1622: data_buf = 8'h16;
			13'h1623: data_buf = 8'h32;
			13'h1624: data_buf = 8'h5a;
			13'h1625: data_buf = 8'h80;
			13'h1626: data_buf = 8'hf1;
			13'h1627: data_buf = 8'hf1;
			13'h1628: data_buf = 8'h37;
			13'h1629: data_buf = 8'hd2;
			13'h162a: data_buf = 8'hc1;
			13'h162b: data_buf = 8'he1;
			13'h162c: data_buf = 8'h79;
			13'h162d: data_buf = 8'h3c;
			13'h162e: data_buf = 8'h3d;
			13'h162f: data_buf = 8'h1f;
			13'h1630: data_buf = 8'hfa;
			13'h1631: data_buf = 8'hdd;
			13'h1632: data_buf = 8'h14;
			13'h1633: data_buf = 8'h17;
			13'h1634: data_buf = 8'h7b;
			13'h1635: data_buf = 8'h17;
			13'h1636: data_buf = 8'h5f;
			13'h1637: data_buf = 8'h7a;
			13'h1638: data_buf = 8'h17;
			13'h1639: data_buf = 8'h57;
			13'h163a: data_buf = 8'h79;
			13'h163b: data_buf = 8'h17;
			13'h163c: data_buf = 8'h4f;
			13'h163d: data_buf = 8'h29;
			13'h163e: data_buf = 8'h78;
			13'h163f: data_buf = 8'h17;
			13'h1640: data_buf = 8'h47;
			13'h1641: data_buf = 8'h3a;
			13'h1642: data_buf = 8'h5a;
			13'h1643: data_buf = 8'h80;
			13'h1644: data_buf = 8'h17;
			13'h1645: data_buf = 8'h32;
			13'h1646: data_buf = 8'h5a;
			13'h1647: data_buf = 8'h80;
			13'h1648: data_buf = 8'h79;
			13'h1649: data_buf = 8'hb2;
			13'h164a: data_buf = 8'hb3;
			13'h164b: data_buf = 8'hc2;
			13'h164c: data_buf = 8'h17;
			13'h164d: data_buf = 8'h16;
			13'h164e: data_buf = 8'he5;
			13'h164f: data_buf = 8'h21;
			13'h1650: data_buf = 8'h2c;
			13'h1651: data_buf = 8'h81;
			13'h1652: data_buf = 8'h35;
			13'h1653: data_buf = 8'he1;
			13'h1654: data_buf = 8'hc2;
			13'h1655: data_buf = 8'h17;
			13'h1656: data_buf = 8'h16;
			13'h1657: data_buf = 8'hc3;
			13'h1658: data_buf = 8'h04;
			13'h1659: data_buf = 8'h04;
			13'h165a: data_buf = 8'h78;
			13'h165b: data_buf = 8'hb7;
			13'h165c: data_buf = 8'hca;
			13'h165d: data_buf = 8'h7e;
			13'h165e: data_buf = 8'h16;
			13'h165f: data_buf = 8'h7d;
			13'h1660: data_buf = 8'h21;
			13'h1661: data_buf = 8'h2c;
			13'h1662: data_buf = 8'h81;
			13'h1663: data_buf = 8'hae;
			13'h1664: data_buf = 8'h80;
			13'h1665: data_buf = 8'h47;
			13'h1666: data_buf = 8'h1f;
			13'h1667: data_buf = 8'ha8;
			13'h1668: data_buf = 8'h78;
			13'h1669: data_buf = 8'hf2;
			13'h166a: data_buf = 8'h7d;
			13'h166b: data_buf = 8'h16;
			13'h166c: data_buf = 8'hc6;
			13'h166d: data_buf = 8'h80;
			13'h166e: data_buf = 8'h77;
			13'h166f: data_buf = 8'hca;
			13'h1670: data_buf = 8'hdd;
			13'h1671: data_buf = 8'h15;
			13'h1672: data_buf = 8'hcd;
			13'h1673: data_buf = 8'h02;
			13'h1674: data_buf = 8'h17;
			13'h1675: data_buf = 8'h77;
			13'h1676: data_buf = 8'h2b;
			13'h1677: data_buf = 8'hc9;
			13'h1678: data_buf = 8'hcd;
			13'h1679: data_buf = 8'h9c;
			13'h167a: data_buf = 8'h16;
			13'h167b: data_buf = 8'h2f;
			13'h167c: data_buf = 8'he1;
			13'h167d: data_buf = 8'hb7;
			13'h167e: data_buf = 8'he1;
			13'h167f: data_buf = 8'hf2;
			13'h1680: data_buf = 8'hbc;
			13'h1681: data_buf = 8'h14;
			13'h1682: data_buf = 8'hc3;
			13'h1683: data_buf = 8'h04;
			13'h1684: data_buf = 8'h04;
			13'h1685: data_buf = 8'hcd;
			13'h1686: data_buf = 8'he8;
			13'h1687: data_buf = 8'h16;
			13'h1688: data_buf = 8'h78;
			13'h1689: data_buf = 8'hb7;
			13'h168a: data_buf = 8'hc8;
			13'h168b: data_buf = 8'hc6;
			13'h168c: data_buf = 8'h02;
			13'h168d: data_buf = 8'hda;
			13'h168e: data_buf = 8'h04;
			13'h168f: data_buf = 8'h04;
			13'h1690: data_buf = 8'h47;
			13'h1691: data_buf = 8'hcd;
			13'h1692: data_buf = 8'h56;
			13'h1693: data_buf = 8'h14;
			13'h1694: data_buf = 8'h21;
			13'h1695: data_buf = 8'h2c;
			13'h1696: data_buf = 8'h81;
			13'h1697: data_buf = 8'h34;
			13'h1698: data_buf = 8'hc0;
			13'h1699: data_buf = 8'hc3;
			13'h169a: data_buf = 8'h04;
			13'h169b: data_buf = 8'h04;
			13'h169c: data_buf = 8'h3a;
			13'h169d: data_buf = 8'h2c;
			13'h169e: data_buf = 8'h81;
			13'h169f: data_buf = 8'hb7;
			13'h16a0: data_buf = 8'hc8;
			13'h16a1: data_buf = 8'h3a;
			13'h16a2: data_buf = 8'h2b;
			13'h16a3: data_buf = 8'h81;
			13'h16a4: data_buf = 8'hfe;
			13'h16a5: data_buf = 8'h2f;
			13'h16a6: data_buf = 8'h17;
			13'h16a7: data_buf = 8'h9f;
			13'h16a8: data_buf = 8'hc0;
			13'h16a9: data_buf = 8'h3c;
			13'h16aa: data_buf = 8'hc9;
			13'h16ab: data_buf = 8'hcd;
			13'h16ac: data_buf = 8'h9c;
			13'h16ad: data_buf = 8'h16;
			13'h16ae: data_buf = 8'h06;
			13'h16af: data_buf = 8'h88;
			13'h16b0: data_buf = 8'h11;
			13'h16b1: data_buf = 8'h00;
			13'h16b2: data_buf = 8'h00;
			13'h16b3: data_buf = 8'h21;
			13'h16b4: data_buf = 8'h2c;
			13'h16b5: data_buf = 8'h81;
			13'h16b6: data_buf = 8'h4f;
			13'h16b7: data_buf = 8'h70;
			13'h16b8: data_buf = 8'h06;
			13'h16b9: data_buf = 8'h00;
			13'h16ba: data_buf = 8'h23;
			13'h16bb: data_buf = 8'h36;
			13'h16bc: data_buf = 8'h80;
			13'h16bd: data_buf = 8'h17;
			13'h16be: data_buf = 8'hc3;
			13'h16bf: data_buf = 8'ha4;
			13'h16c0: data_buf = 8'h14;
			13'h16c1: data_buf = 8'hcd;
			13'h16c2: data_buf = 8'h9c;
			13'h16c3: data_buf = 8'h16;
			13'h16c4: data_buf = 8'hf0;
			13'h16c5: data_buf = 8'h21;
			13'h16c6: data_buf = 8'h2b;
			13'h16c7: data_buf = 8'h81;
			13'h16c8: data_buf = 8'h7e;
			13'h16c9: data_buf = 8'hee;
			13'h16ca: data_buf = 8'h80;
			13'h16cb: data_buf = 8'h77;
			13'h16cc: data_buf = 8'hc9;
			13'h16cd: data_buf = 8'heb;
			13'h16ce: data_buf = 8'h2a;
			13'h16cf: data_buf = 8'h29;
			13'h16d0: data_buf = 8'h81;
			13'h16d1: data_buf = 8'he3;
			13'h16d2: data_buf = 8'he5;
			13'h16d3: data_buf = 8'h2a;
			13'h16d4: data_buf = 8'h2b;
			13'h16d5: data_buf = 8'h81;
			13'h16d6: data_buf = 8'he3;
			13'h16d7: data_buf = 8'he5;
			13'h16d8: data_buf = 8'heb;
			13'h16d9: data_buf = 8'hc9;
			13'h16da: data_buf = 8'hcd;
			13'h16db: data_buf = 8'heb;
			13'h16dc: data_buf = 8'h16;
			13'h16dd: data_buf = 8'heb;
			13'h16de: data_buf = 8'h22;
			13'h16df: data_buf = 8'h29;
			13'h16e0: data_buf = 8'h81;
			13'h16e1: data_buf = 8'h60;
			13'h16e2: data_buf = 8'h69;
			13'h16e3: data_buf = 8'h22;
			13'h16e4: data_buf = 8'h2b;
			13'h16e5: data_buf = 8'h81;
			13'h16e6: data_buf = 8'heb;
			13'h16e7: data_buf = 8'hc9;
			13'h16e8: data_buf = 8'h21;
			13'h16e9: data_buf = 8'h29;
			13'h16ea: data_buf = 8'h81;
			13'h16eb: data_buf = 8'h5e;
			13'h16ec: data_buf = 8'h23;
			13'h16ed: data_buf = 8'h56;
			13'h16ee: data_buf = 8'h23;
			13'h16ef: data_buf = 8'h4e;
			13'h16f0: data_buf = 8'h23;
			13'h16f1: data_buf = 8'h46;
			13'h16f2: data_buf = 8'h23;
			13'h16f3: data_buf = 8'hc9;
			13'h16f4: data_buf = 8'h11;
			13'h16f5: data_buf = 8'h29;
			13'h16f6: data_buf = 8'h81;
			13'h16f7: data_buf = 8'h06;
			13'h16f8: data_buf = 8'h04;
			13'h16f9: data_buf = 8'h1a;
			13'h16fa: data_buf = 8'h77;
			13'h16fb: data_buf = 8'h13;
			13'h16fc: data_buf = 8'h23;
			13'h16fd: data_buf = 8'h05;
			13'h16fe: data_buf = 8'hc2;
			13'h16ff: data_buf = 8'hf9;
			13'h1700: data_buf = 8'h16;
			13'h1701: data_buf = 8'hc9;
			13'h1702: data_buf = 8'h21;
			13'h1703: data_buf = 8'h2b;
			13'h1704: data_buf = 8'h81;
			13'h1705: data_buf = 8'h7e;
			13'h1706: data_buf = 8'h07;
			13'h1707: data_buf = 8'h37;
			13'h1708: data_buf = 8'h1f;
			13'h1709: data_buf = 8'h77;
			13'h170a: data_buf = 8'h3f;
			13'h170b: data_buf = 8'h1f;
			13'h170c: data_buf = 8'h23;
			13'h170d: data_buf = 8'h23;
			13'h170e: data_buf = 8'h77;
			13'h170f: data_buf = 8'h79;
			13'h1710: data_buf = 8'h07;
			13'h1711: data_buf = 8'h37;
			13'h1712: data_buf = 8'h1f;
			13'h1713: data_buf = 8'h4f;
			13'h1714: data_buf = 8'h1f;
			13'h1715: data_buf = 8'hae;
			13'h1716: data_buf = 8'hc9;
			13'h1717: data_buf = 8'h78;
			13'h1718: data_buf = 8'hb7;
			13'h1719: data_buf = 8'hca;
			13'h171a: data_buf = 8'h9c;
			13'h171b: data_buf = 8'h16;
			13'h171c: data_buf = 8'h21;
			13'h171d: data_buf = 8'ha5;
			13'h171e: data_buf = 8'h16;
			13'h171f: data_buf = 8'he5;
			13'h1720: data_buf = 8'hcd;
			13'h1721: data_buf = 8'h9c;
			13'h1722: data_buf = 8'h16;
			13'h1723: data_buf = 8'h79;
			13'h1724: data_buf = 8'hc8;
			13'h1725: data_buf = 8'h21;
			13'h1726: data_buf = 8'h2b;
			13'h1727: data_buf = 8'h81;
			13'h1728: data_buf = 8'hae;
			13'h1729: data_buf = 8'h79;
			13'h172a: data_buf = 8'hf8;
			13'h172b: data_buf = 8'hcd;
			13'h172c: data_buf = 8'h31;
			13'h172d: data_buf = 8'h17;
			13'h172e: data_buf = 8'h1f;
			13'h172f: data_buf = 8'ha9;
			13'h1730: data_buf = 8'hc9;
			13'h1731: data_buf = 8'h23;
			13'h1732: data_buf = 8'h78;
			13'h1733: data_buf = 8'hbe;
			13'h1734: data_buf = 8'hc0;
			13'h1735: data_buf = 8'h2b;
			13'h1736: data_buf = 8'h79;
			13'h1737: data_buf = 8'hbe;
			13'h1738: data_buf = 8'hc0;
			13'h1739: data_buf = 8'h2b;
			13'h173a: data_buf = 8'h7a;
			13'h173b: data_buf = 8'hbe;
			13'h173c: data_buf = 8'hc0;
			13'h173d: data_buf = 8'h2b;
			13'h173e: data_buf = 8'h7b;
			13'h173f: data_buf = 8'h96;
			13'h1740: data_buf = 8'hc0;
			13'h1741: data_buf = 8'he1;
			13'h1742: data_buf = 8'he1;
			13'h1743: data_buf = 8'hc9;
			13'h1744: data_buf = 8'h47;
			13'h1745: data_buf = 8'h4f;
			13'h1746: data_buf = 8'h57;
			13'h1747: data_buf = 8'h5f;
			13'h1748: data_buf = 8'hb7;
			13'h1749: data_buf = 8'hc8;
			13'h174a: data_buf = 8'he5;
			13'h174b: data_buf = 8'hcd;
			13'h174c: data_buf = 8'he8;
			13'h174d: data_buf = 8'h16;
			13'h174e: data_buf = 8'hcd;
			13'h174f: data_buf = 8'h02;
			13'h1750: data_buf = 8'h17;
			13'h1751: data_buf = 8'hae;
			13'h1752: data_buf = 8'h67;
			13'h1753: data_buf = 8'hfc;
			13'h1754: data_buf = 8'h68;
			13'h1755: data_buf = 8'h17;
			13'h1756: data_buf = 8'h3e;
			13'h1757: data_buf = 8'h98;
			13'h1758: data_buf = 8'h90;
			13'h1759: data_buf = 8'hcd;
			13'h175a: data_buf = 8'h1b;
			13'h175b: data_buf = 8'h15;
			13'h175c: data_buf = 8'h7c;
			13'h175d: data_buf = 8'h17;
			13'h175e: data_buf = 8'hdc;
			13'h175f: data_buf = 8'hee;
			13'h1760: data_buf = 8'h14;
			13'h1761: data_buf = 8'h06;
			13'h1762: data_buf = 8'h00;
			13'h1763: data_buf = 8'hdc;
			13'h1764: data_buf = 8'h07;
			13'h1765: data_buf = 8'h15;
			13'h1766: data_buf = 8'he1;
			13'h1767: data_buf = 8'hc9;
			13'h1768: data_buf = 8'h1b;
			13'h1769: data_buf = 8'h7a;
			13'h176a: data_buf = 8'ha3;
			13'h176b: data_buf = 8'h3c;
			13'h176c: data_buf = 8'hc0;
			13'h176d: data_buf = 8'h0b;
			13'h176e: data_buf = 8'hc9;
			13'h176f: data_buf = 8'h21;
			13'h1770: data_buf = 8'h2c;
			13'h1771: data_buf = 8'h81;
			13'h1772: data_buf = 8'h7e;
			13'h1773: data_buf = 8'hfe;
			13'h1774: data_buf = 8'h98;
			13'h1775: data_buf = 8'h3a;
			13'h1776: data_buf = 8'h29;
			13'h1777: data_buf = 8'h81;
			13'h1778: data_buf = 8'hd0;
			13'h1779: data_buf = 8'h7e;
			13'h177a: data_buf = 8'hcd;
			13'h177b: data_buf = 8'h44;
			13'h177c: data_buf = 8'h17;
			13'h177d: data_buf = 8'h36;
			13'h177e: data_buf = 8'h98;
			13'h177f: data_buf = 8'h7b;
			13'h1780: data_buf = 8'hf5;
			13'h1781: data_buf = 8'h79;
			13'h1782: data_buf = 8'h17;
			13'h1783: data_buf = 8'hcd;
			13'h1784: data_buf = 8'ha4;
			13'h1785: data_buf = 8'h14;
			13'h1786: data_buf = 8'hf1;
			13'h1787: data_buf = 8'hc9;
			13'h1788: data_buf = 8'h21;
			13'h1789: data_buf = 8'h00;
			13'h178a: data_buf = 8'h00;
			13'h178b: data_buf = 8'h78;
			13'h178c: data_buf = 8'hb1;
			13'h178d: data_buf = 8'hc8;
			13'h178e: data_buf = 8'h3e;
			13'h178f: data_buf = 8'h10;
			13'h1790: data_buf = 8'h29;
			13'h1791: data_buf = 8'hda;
			13'h1792: data_buf = 8'hc8;
			13'h1793: data_buf = 8'h0f;
			13'h1794: data_buf = 8'heb;
			13'h1795: data_buf = 8'h29;
			13'h1796: data_buf = 8'heb;
			13'h1797: data_buf = 8'hd2;
			13'h1798: data_buf = 8'h9e;
			13'h1799: data_buf = 8'h17;
			13'h179a: data_buf = 8'h09;
			13'h179b: data_buf = 8'hda;
			13'h179c: data_buf = 8'hc8;
			13'h179d: data_buf = 8'h0f;
			13'h179e: data_buf = 8'h3d;
			13'h179f: data_buf = 8'hc2;
			13'h17a0: data_buf = 8'h90;
			13'h17a1: data_buf = 8'h17;
			13'h17a2: data_buf = 8'hc9;
			13'h17a3: data_buf = 8'hfe;
			13'h17a4: data_buf = 8'h2d;
			13'h17a5: data_buf = 8'hf5;
			13'h17a6: data_buf = 8'hca;
			13'h17a7: data_buf = 8'haf;
			13'h17a8: data_buf = 8'h17;
			13'h17a9: data_buf = 8'hfe;
			13'h17aa: data_buf = 8'h2b;
			13'h17ab: data_buf = 8'hca;
			13'h17ac: data_buf = 8'haf;
			13'h17ad: data_buf = 8'h17;
			13'h17ae: data_buf = 8'h2b;
			13'h17af: data_buf = 8'hcd;
			13'h17b0: data_buf = 8'hbc;
			13'h17b1: data_buf = 8'h14;
			13'h17b2: data_buf = 8'h47;
			13'h17b3: data_buf = 8'h57;
			13'h17b4: data_buf = 8'h5f;
			13'h17b5: data_buf = 8'h2f;
			13'h17b6: data_buf = 8'h4f;
			13'h17b7: data_buf = 8'hcd;
			13'h17b8: data_buf = 8'h4d;
			13'h17b9: data_buf = 8'h08;
			13'h17ba: data_buf = 8'hda;
			13'h17bb: data_buf = 8'h00;
			13'h17bc: data_buf = 8'h18;
			13'h17bd: data_buf = 8'hfe;
			13'h17be: data_buf = 8'h2e;
			13'h17bf: data_buf = 8'hca;
			13'h17c0: data_buf = 8'hdb;
			13'h17c1: data_buf = 8'h17;
			13'h17c2: data_buf = 8'hfe;
			13'h17c3: data_buf = 8'h45;
			13'h17c4: data_buf = 8'hc2;
			13'h17c5: data_buf = 8'hdf;
			13'h17c6: data_buf = 8'h17;
			13'h17c7: data_buf = 8'hcd;
			13'h17c8: data_buf = 8'h4d;
			13'h17c9: data_buf = 8'h08;
			13'h17ca: data_buf = 8'hcd;
			13'h17cb: data_buf = 8'hf3;
			13'h17cc: data_buf = 8'h0d;
			13'h17cd: data_buf = 8'hcd;
			13'h17ce: data_buf = 8'h4d;
			13'h17cf: data_buf = 8'h08;
			13'h17d0: data_buf = 8'hda;
			13'h17d1: data_buf = 8'h22;
			13'h17d2: data_buf = 8'h18;
			13'h17d3: data_buf = 8'h14;
			13'h17d4: data_buf = 8'hc2;
			13'h17d5: data_buf = 8'hdf;
			13'h17d6: data_buf = 8'h17;
			13'h17d7: data_buf = 8'haf;
			13'h17d8: data_buf = 8'h93;
			13'h17d9: data_buf = 8'h5f;
			13'h17da: data_buf = 8'h0c;
			13'h17db: data_buf = 8'h0c;
			13'h17dc: data_buf = 8'hca;
			13'h17dd: data_buf = 8'hb7;
			13'h17de: data_buf = 8'h17;
			13'h17df: data_buf = 8'he5;
			13'h17e0: data_buf = 8'h7b;
			13'h17e1: data_buf = 8'h90;
			13'h17e2: data_buf = 8'hf4;
			13'h17e3: data_buf = 8'hf8;
			13'h17e4: data_buf = 8'h17;
			13'h17e5: data_buf = 8'hf2;
			13'h17e6: data_buf = 8'hee;
			13'h17e7: data_buf = 8'h17;
			13'h17e8: data_buf = 8'hf5;
			13'h17e9: data_buf = 8'hcd;
			13'h17ea: data_buf = 8'he4;
			13'h17eb: data_buf = 8'h15;
			13'h17ec: data_buf = 8'hf1;
			13'h17ed: data_buf = 8'h3c;
			13'h17ee: data_buf = 8'hc2;
			13'h17ef: data_buf = 8'he2;
			13'h17f0: data_buf = 8'h17;
			13'h17f1: data_buf = 8'hd1;
			13'h17f2: data_buf = 8'hf1;
			13'h17f3: data_buf = 8'hcc;
			13'h17f4: data_buf = 8'hc5;
			13'h17f5: data_buf = 8'h16;
			13'h17f6: data_buf = 8'heb;
			13'h17f7: data_buf = 8'hc9;
			13'h17f8: data_buf = 8'hc8;
			13'h17f9: data_buf = 8'hf5;
			13'h17fa: data_buf = 8'hcd;
			13'h17fb: data_buf = 8'h85;
			13'h17fc: data_buf = 8'h16;
			13'h17fd: data_buf = 8'hf1;
			13'h17fe: data_buf = 8'h3d;
			13'h17ff: data_buf = 8'hc9;
			13'h1800: data_buf = 8'hd5;
			13'h1801: data_buf = 8'h57;
			13'h1802: data_buf = 8'h78;
			13'h1803: data_buf = 8'h89;
			13'h1804: data_buf = 8'h47;
			13'h1805: data_buf = 8'hc5;
			13'h1806: data_buf = 8'he5;
			13'h1807: data_buf = 8'hd5;
			13'h1808: data_buf = 8'hcd;
			13'h1809: data_buf = 8'h85;
			13'h180a: data_buf = 8'h16;
			13'h180b: data_buf = 8'hf1;
			13'h180c: data_buf = 8'hd6;
			13'h180d: data_buf = 8'h30;
			13'h180e: data_buf = 8'hcd;
			13'h180f: data_buf = 8'h17;
			13'h1810: data_buf = 8'h18;
			13'h1811: data_buf = 8'he1;
			13'h1812: data_buf = 8'hc1;
			13'h1813: data_buf = 8'hd1;
			13'h1814: data_buf = 8'hc3;
			13'h1815: data_buf = 8'hb7;
			13'h1816: data_buf = 8'h17;
			13'h1817: data_buf = 8'hcd;
			13'h1818: data_buf = 8'hcd;
			13'h1819: data_buf = 8'h16;
			13'h181a: data_buf = 8'hcd;
			13'h181b: data_buf = 8'hae;
			13'h181c: data_buf = 8'h16;
			13'h181d: data_buf = 8'hc1;
			13'h181e: data_buf = 8'hd1;
			13'h181f: data_buf = 8'hc3;
			13'h1820: data_buf = 8'h56;
			13'h1821: data_buf = 8'h14;
			13'h1822: data_buf = 8'h7b;
			13'h1823: data_buf = 8'h07;
			13'h1824: data_buf = 8'h07;
			13'h1825: data_buf = 8'h83;
			13'h1826: data_buf = 8'h07;
			13'h1827: data_buf = 8'h86;
			13'h1828: data_buf = 8'hd6;
			13'h1829: data_buf = 8'h30;
			13'h182a: data_buf = 8'h5f;
			13'h182b: data_buf = 8'hc3;
			13'h182c: data_buf = 8'hcd;
			13'h182d: data_buf = 8'h17;
			13'h182e: data_buf = 8'he5;
			13'h182f: data_buf = 8'h21;
			13'h1830: data_buf = 8'h8d;
			13'h1831: data_buf = 8'h03;
			13'h1832: data_buf = 8'hcd;
			13'h1833: data_buf = 8'h93;
			13'h1834: data_buf = 8'h11;
			13'h1835: data_buf = 8'he1;
			13'h1836: data_buf = 8'heb;
			13'h1837: data_buf = 8'haf;
			13'h1838: data_buf = 8'h06;
			13'h1839: data_buf = 8'h98;
			13'h183a: data_buf = 8'hcd;
			13'h183b: data_buf = 8'hb3;
			13'h183c: data_buf = 8'h16;
			13'h183d: data_buf = 8'h21;
			13'h183e: data_buf = 8'h92;
			13'h183f: data_buf = 8'h11;
			13'h1840: data_buf = 8'he5;
			13'h1841: data_buf = 8'h21;
			13'h1842: data_buf = 8'h2e;
			13'h1843: data_buf = 8'h81;
			13'h1844: data_buf = 8'he5;
			13'h1845: data_buf = 8'hcd;
			13'h1846: data_buf = 8'h9c;
			13'h1847: data_buf = 8'h16;
			13'h1848: data_buf = 8'h36;
			13'h1849: data_buf = 8'h20;
			13'h184a: data_buf = 8'hf2;
			13'h184b: data_buf = 8'h4f;
			13'h184c: data_buf = 8'h18;
			13'h184d: data_buf = 8'h36;
			13'h184e: data_buf = 8'h2d;
			13'h184f: data_buf = 8'h23;
			13'h1850: data_buf = 8'h36;
			13'h1851: data_buf = 8'h30;
			13'h1852: data_buf = 8'hca;
			13'h1853: data_buf = 8'h05;
			13'h1854: data_buf = 8'h19;
			13'h1855: data_buf = 8'he5;
			13'h1856: data_buf = 8'hfc;
			13'h1857: data_buf = 8'hc5;
			13'h1858: data_buf = 8'h16;
			13'h1859: data_buf = 8'haf;
			13'h185a: data_buf = 8'hf5;
			13'h185b: data_buf = 8'hcd;
			13'h185c: data_buf = 8'h0b;
			13'h185d: data_buf = 8'h19;
			13'h185e: data_buf = 8'h01;
			13'h185f: data_buf = 8'h43;
			13'h1860: data_buf = 8'h91;
			13'h1861: data_buf = 8'h11;
			13'h1862: data_buf = 8'hf8;
			13'h1863: data_buf = 8'h4f;
			13'h1864: data_buf = 8'hcd;
			13'h1865: data_buf = 8'h17;
			13'h1866: data_buf = 8'h17;
			13'h1867: data_buf = 8'hb7;
			13'h1868: data_buf = 8'he2;
			13'h1869: data_buf = 8'h7c;
			13'h186a: data_buf = 8'h18;
			13'h186b: data_buf = 8'hf1;
			13'h186c: data_buf = 8'hcd;
			13'h186d: data_buf = 8'hf9;
			13'h186e: data_buf = 8'h17;
			13'h186f: data_buf = 8'hf5;
			13'h1870: data_buf = 8'hc3;
			13'h1871: data_buf = 8'h5e;
			13'h1872: data_buf = 8'h18;
			13'h1873: data_buf = 8'hcd;
			13'h1874: data_buf = 8'he4;
			13'h1875: data_buf = 8'h15;
			13'h1876: data_buf = 8'hf1;
			13'h1877: data_buf = 8'h3c;
			13'h1878: data_buf = 8'hf5;
			13'h1879: data_buf = 8'hcd;
			13'h187a: data_buf = 8'h0b;
			13'h187b: data_buf = 8'h19;
			13'h187c: data_buf = 8'hcd;
			13'h187d: data_buf = 8'h44;
			13'h187e: data_buf = 8'h14;
			13'h187f: data_buf = 8'h3c;
			13'h1880: data_buf = 8'hcd;
			13'h1881: data_buf = 8'h44;
			13'h1882: data_buf = 8'h17;
			13'h1883: data_buf = 8'hcd;
			13'h1884: data_buf = 8'hdd;
			13'h1885: data_buf = 8'h16;
			13'h1886: data_buf = 8'h01;
			13'h1887: data_buf = 8'h06;
			13'h1888: data_buf = 8'h03;
			13'h1889: data_buf = 8'hf1;
			13'h188a: data_buf = 8'h81;
			13'h188b: data_buf = 8'h3c;
			13'h188c: data_buf = 8'hfa;
			13'h188d: data_buf = 8'h98;
			13'h188e: data_buf = 8'h18;
			13'h188f: data_buf = 8'hfe;
			13'h1890: data_buf = 8'h08;
			13'h1891: data_buf = 8'hd2;
			13'h1892: data_buf = 8'h98;
			13'h1893: data_buf = 8'h18;
			13'h1894: data_buf = 8'h3c;
			13'h1895: data_buf = 8'h47;
			13'h1896: data_buf = 8'h3e;
			13'h1897: data_buf = 8'h02;
			13'h1898: data_buf = 8'h3d;
			13'h1899: data_buf = 8'h3d;
			13'h189a: data_buf = 8'he1;
			13'h189b: data_buf = 8'hf5;
			13'h189c: data_buf = 8'h11;
			13'h189d: data_buf = 8'h1e;
			13'h189e: data_buf = 8'h19;
			13'h189f: data_buf = 8'h05;
			13'h18a0: data_buf = 8'hc2;
			13'h18a1: data_buf = 8'ha9;
			13'h18a2: data_buf = 8'h18;
			13'h18a3: data_buf = 8'h36;
			13'h18a4: data_buf = 8'h2e;
			13'h18a5: data_buf = 8'h23;
			13'h18a6: data_buf = 8'h36;
			13'h18a7: data_buf = 8'h30;
			13'h18a8: data_buf = 8'h23;
			13'h18a9: data_buf = 8'h05;
			13'h18aa: data_buf = 8'h36;
			13'h18ab: data_buf = 8'h2e;
			13'h18ac: data_buf = 8'hcc;
			13'h18ad: data_buf = 8'hf2;
			13'h18ae: data_buf = 8'h16;
			13'h18af: data_buf = 8'hc5;
			13'h18b0: data_buf = 8'he5;
			13'h18b1: data_buf = 8'hd5;
			13'h18b2: data_buf = 8'hcd;
			13'h18b3: data_buf = 8'he8;
			13'h18b4: data_buf = 8'h16;
			13'h18b5: data_buf = 8'he1;
			13'h18b6: data_buf = 8'h06;
			13'h18b7: data_buf = 8'h2f;
			13'h18b8: data_buf = 8'h04;
			13'h18b9: data_buf = 8'h7b;
			13'h18ba: data_buf = 8'h96;
			13'h18bb: data_buf = 8'h5f;
			13'h18bc: data_buf = 8'h23;
			13'h18bd: data_buf = 8'h7a;
			13'h18be: data_buf = 8'h9e;
			13'h18bf: data_buf = 8'h57;
			13'h18c0: data_buf = 8'h23;
			13'h18c1: data_buf = 8'h79;
			13'h18c2: data_buf = 8'h9e;
			13'h18c3: data_buf = 8'h4f;
			13'h18c4: data_buf = 8'h2b;
			13'h18c5: data_buf = 8'h2b;
			13'h18c6: data_buf = 8'hd2;
			13'h18c7: data_buf = 8'hb8;
			13'h18c8: data_buf = 8'h18;
			13'h18c9: data_buf = 8'hcd;
			13'h18ca: data_buf = 8'hfb;
			13'h18cb: data_buf = 8'h14;
			13'h18cc: data_buf = 8'h23;
			13'h18cd: data_buf = 8'hcd;
			13'h18ce: data_buf = 8'hdd;
			13'h18cf: data_buf = 8'h16;
			13'h18d0: data_buf = 8'heb;
			13'h18d1: data_buf = 8'he1;
			13'h18d2: data_buf = 8'h70;
			13'h18d3: data_buf = 8'h23;
			13'h18d4: data_buf = 8'hc1;
			13'h18d5: data_buf = 8'h0d;
			13'h18d6: data_buf = 8'hc2;
			13'h18d7: data_buf = 8'ha9;
			13'h18d8: data_buf = 8'h18;
			13'h18d9: data_buf = 8'h05;
			13'h18da: data_buf = 8'hca;
			13'h18db: data_buf = 8'he9;
			13'h18dc: data_buf = 8'h18;
			13'h18dd: data_buf = 8'h2b;
			13'h18de: data_buf = 8'h7e;
			13'h18df: data_buf = 8'hfe;
			13'h18e0: data_buf = 8'h30;
			13'h18e1: data_buf = 8'hca;
			13'h18e2: data_buf = 8'hdd;
			13'h18e3: data_buf = 8'h18;
			13'h18e4: data_buf = 8'hfe;
			13'h18e5: data_buf = 8'h2e;
			13'h18e6: data_buf = 8'hc4;
			13'h18e7: data_buf = 8'hf2;
			13'h18e8: data_buf = 8'h16;
			13'h18e9: data_buf = 8'hf1;
			13'h18ea: data_buf = 8'hca;
			13'h18eb: data_buf = 8'h08;
			13'h18ec: data_buf = 8'h19;
			13'h18ed: data_buf = 8'h36;
			13'h18ee: data_buf = 8'h45;
			13'h18ef: data_buf = 8'h23;
			13'h18f0: data_buf = 8'h36;
			13'h18f1: data_buf = 8'h2b;
			13'h18f2: data_buf = 8'hf2;
			13'h18f3: data_buf = 8'hf9;
			13'h18f4: data_buf = 8'h18;
			13'h18f5: data_buf = 8'h36;
			13'h18f6: data_buf = 8'h2d;
			13'h18f7: data_buf = 8'h2f;
			13'h18f8: data_buf = 8'h3c;
			13'h18f9: data_buf = 8'h06;
			13'h18fa: data_buf = 8'h2f;
			13'h18fb: data_buf = 8'h04;
			13'h18fc: data_buf = 8'hd6;
			13'h18fd: data_buf = 8'h0a;
			13'h18fe: data_buf = 8'hd2;
			13'h18ff: data_buf = 8'hfb;
			13'h1900: data_buf = 8'h18;
			13'h1901: data_buf = 8'hc6;
			13'h1902: data_buf = 8'h3a;
			13'h1903: data_buf = 8'h23;
			13'h1904: data_buf = 8'h70;
			13'h1905: data_buf = 8'h23;
			13'h1906: data_buf = 8'h77;
			13'h1907: data_buf = 8'h23;
			13'h1908: data_buf = 8'h71;
			13'h1909: data_buf = 8'he1;
			13'h190a: data_buf = 8'hc9;
			13'h190b: data_buf = 8'h01;
			13'h190c: data_buf = 8'h74;
			13'h190d: data_buf = 8'h94;
			13'h190e: data_buf = 8'h11;
			13'h190f: data_buf = 8'hf7;
			13'h1910: data_buf = 8'h23;
			13'h1911: data_buf = 8'hcd;
			13'h1912: data_buf = 8'h17;
			13'h1913: data_buf = 8'h17;
			13'h1914: data_buf = 8'hb7;
			13'h1915: data_buf = 8'he1;
			13'h1916: data_buf = 8'he2;
			13'h1917: data_buf = 8'h73;
			13'h1918: data_buf = 8'h18;
			13'h1919: data_buf = 8'he9;
			13'h191a: data_buf = 8'h00;
			13'h191b: data_buf = 8'h00;
			13'h191c: data_buf = 8'h00;
			13'h191d: data_buf = 8'h80;
			13'h191e: data_buf = 8'ha0;
			13'h191f: data_buf = 8'h86;
			13'h1920: data_buf = 8'h01;
			13'h1921: data_buf = 8'h10;
			13'h1922: data_buf = 8'h27;
			13'h1923: data_buf = 8'h00;
			13'h1924: data_buf = 8'he8;
			13'h1925: data_buf = 8'h03;
			13'h1926: data_buf = 8'h00;
			13'h1927: data_buf = 8'h64;
			13'h1928: data_buf = 8'h00;
			13'h1929: data_buf = 8'h00;
			13'h192a: data_buf = 8'h0a;
			13'h192b: data_buf = 8'h00;
			13'h192c: data_buf = 8'h00;
			13'h192d: data_buf = 8'h01;
			13'h192e: data_buf = 8'h00;
			13'h192f: data_buf = 8'h00;
			13'h1930: data_buf = 8'h21;
			13'h1931: data_buf = 8'hc5;
			13'h1932: data_buf = 8'h16;
			13'h1933: data_buf = 8'he3;
			13'h1934: data_buf = 8'he9;
			13'h1935: data_buf = 8'hcd;
			13'h1936: data_buf = 8'hcd;
			13'h1937: data_buf = 8'h16;
			13'h1938: data_buf = 8'h21;
			13'h1939: data_buf = 8'h1a;
			13'h193a: data_buf = 8'h19;
			13'h193b: data_buf = 8'hcd;
			13'h193c: data_buf = 8'hda;
			13'h193d: data_buf = 8'h16;
			13'h193e: data_buf = 8'hc1;
			13'h193f: data_buf = 8'hd1;
			13'h1940: data_buf = 8'hcd;
			13'h1941: data_buf = 8'h9c;
			13'h1942: data_buf = 8'h16;
			13'h1943: data_buf = 8'h78;
			13'h1944: data_buf = 8'hca;
			13'h1945: data_buf = 8'h83;
			13'h1946: data_buf = 8'h19;
			13'h1947: data_buf = 8'hf2;
			13'h1948: data_buf = 8'h4e;
			13'h1949: data_buf = 8'h19;
			13'h194a: data_buf = 8'hb7;
			13'h194b: data_buf = 8'hca;
			13'h194c: data_buf = 8'hf8;
			13'h194d: data_buf = 8'h03;
			13'h194e: data_buf = 8'hb7;
			13'h194f: data_buf = 8'hca;
			13'h1950: data_buf = 8'hbd;
			13'h1951: data_buf = 8'h14;
			13'h1952: data_buf = 8'hd5;
			13'h1953: data_buf = 8'hc5;
			13'h1954: data_buf = 8'h79;
			13'h1955: data_buf = 8'hf6;
			13'h1956: data_buf = 8'h7f;
			13'h1957: data_buf = 8'hcd;
			13'h1958: data_buf = 8'he8;
			13'h1959: data_buf = 8'h16;
			13'h195a: data_buf = 8'hf2;
			13'h195b: data_buf = 8'h6b;
			13'h195c: data_buf = 8'h19;
			13'h195d: data_buf = 8'hd5;
			13'h195e: data_buf = 8'hc5;
			13'h195f: data_buf = 8'hcd;
			13'h1960: data_buf = 8'h6f;
			13'h1961: data_buf = 8'h17;
			13'h1962: data_buf = 8'hc1;
			13'h1963: data_buf = 8'hd1;
			13'h1964: data_buf = 8'hf5;
			13'h1965: data_buf = 8'hcd;
			13'h1966: data_buf = 8'h17;
			13'h1967: data_buf = 8'h17;
			13'h1968: data_buf = 8'he1;
			13'h1969: data_buf = 8'h7c;
			13'h196a: data_buf = 8'h1f;
			13'h196b: data_buf = 8'he1;
			13'h196c: data_buf = 8'h22;
			13'h196d: data_buf = 8'h2b;
			13'h196e: data_buf = 8'h81;
			13'h196f: data_buf = 8'he1;
			13'h1970: data_buf = 8'h22;
			13'h1971: data_buf = 8'h29;
			13'h1972: data_buf = 8'h81;
			13'h1973: data_buf = 8'hdc;
			13'h1974: data_buf = 8'h30;
			13'h1975: data_buf = 8'h19;
			13'h1976: data_buf = 8'hcc;
			13'h1977: data_buf = 8'hc5;
			13'h1978: data_buf = 8'h16;
			13'h1979: data_buf = 8'hd5;
			13'h197a: data_buf = 8'hc5;
			13'h197b: data_buf = 8'hcd;
			13'h197c: data_buf = 8'h50;
			13'h197d: data_buf = 8'h15;
			13'h197e: data_buf = 8'hc1;
			13'h197f: data_buf = 8'hd1;
			13'h1980: data_buf = 8'hcd;
			13'h1981: data_buf = 8'h91;
			13'h1982: data_buf = 8'h15;
			13'h1983: data_buf = 8'hcd;
			13'h1984: data_buf = 8'hcd;
			13'h1985: data_buf = 8'h16;
			13'h1986: data_buf = 8'h01;
			13'h1987: data_buf = 8'h38;
			13'h1988: data_buf = 8'h81;
			13'h1989: data_buf = 8'h11;
			13'h198a: data_buf = 8'h3b;
			13'h198b: data_buf = 8'haa;
			13'h198c: data_buf = 8'hcd;
			13'h198d: data_buf = 8'h91;
			13'h198e: data_buf = 8'h15;
			13'h198f: data_buf = 8'h3a;
			13'h1990: data_buf = 8'h2c;
			13'h1991: data_buf = 8'h81;
			13'h1992: data_buf = 8'hfe;
			13'h1993: data_buf = 8'h88;
			13'h1994: data_buf = 8'hd2;
			13'h1995: data_buf = 8'h78;
			13'h1996: data_buf = 8'h16;
			13'h1997: data_buf = 8'hcd;
			13'h1998: data_buf = 8'h6f;
			13'h1999: data_buf = 8'h17;
			13'h199a: data_buf = 8'hc6;
			13'h199b: data_buf = 8'h80;
			13'h199c: data_buf = 8'hc6;
			13'h199d: data_buf = 8'h02;
			13'h199e: data_buf = 8'hda;
			13'h199f: data_buf = 8'h78;
			13'h19a0: data_buf = 8'h16;
			13'h19a1: data_buf = 8'hf5;
			13'h19a2: data_buf = 8'h21;
			13'h19a3: data_buf = 8'h3f;
			13'h19a4: data_buf = 8'h15;
			13'h19a5: data_buf = 8'hcd;
			13'h19a6: data_buf = 8'h47;
			13'h19a7: data_buf = 8'h14;
			13'h19a8: data_buf = 8'hcd;
			13'h19a9: data_buf = 8'h88;
			13'h19aa: data_buf = 8'h15;
			13'h19ab: data_buf = 8'hf1;
			13'h19ac: data_buf = 8'hc1;
			13'h19ad: data_buf = 8'hd1;
			13'h19ae: data_buf = 8'hf5;
			13'h19af: data_buf = 8'hcd;
			13'h19b0: data_buf = 8'h53;
			13'h19b1: data_buf = 8'h14;
			13'h19b2: data_buf = 8'hcd;
			13'h19b3: data_buf = 8'hc5;
			13'h19b4: data_buf = 8'h16;
			13'h19b5: data_buf = 8'h21;
			13'h19b6: data_buf = 8'hc3;
			13'h19b7: data_buf = 8'h19;
			13'h19b8: data_buf = 8'hcd;
			13'h19b9: data_buf = 8'hf3;
			13'h19ba: data_buf = 8'h19;
			13'h19bb: data_buf = 8'h11;
			13'h19bc: data_buf = 8'h00;
			13'h19bd: data_buf = 8'h00;
			13'h19be: data_buf = 8'hc1;
			13'h19bf: data_buf = 8'h4a;
			13'h19c0: data_buf = 8'hc3;
			13'h19c1: data_buf = 8'h91;
			13'h19c2: data_buf = 8'h15;
			13'h19c3: data_buf = 8'h08;
			13'h19c4: data_buf = 8'h40;
			13'h19c5: data_buf = 8'h2e;
			13'h19c6: data_buf = 8'h94;
			13'h19c7: data_buf = 8'h74;
			13'h19c8: data_buf = 8'h70;
			13'h19c9: data_buf = 8'h4f;
			13'h19ca: data_buf = 8'h2e;
			13'h19cb: data_buf = 8'h77;
			13'h19cc: data_buf = 8'h6e;
			13'h19cd: data_buf = 8'h02;
			13'h19ce: data_buf = 8'h88;
			13'h19cf: data_buf = 8'h7a;
			13'h19d0: data_buf = 8'he6;
			13'h19d1: data_buf = 8'ha0;
			13'h19d2: data_buf = 8'h2a;
			13'h19d3: data_buf = 8'h7c;
			13'h19d4: data_buf = 8'h50;
			13'h19d5: data_buf = 8'haa;
			13'h19d6: data_buf = 8'haa;
			13'h19d7: data_buf = 8'h7e;
			13'h19d8: data_buf = 8'hff;
			13'h19d9: data_buf = 8'hff;
			13'h19da: data_buf = 8'h7f;
			13'h19db: data_buf = 8'h7f;
			13'h19dc: data_buf = 8'h00;
			13'h19dd: data_buf = 8'h00;
			13'h19de: data_buf = 8'h80;
			13'h19df: data_buf = 8'h81;
			13'h19e0: data_buf = 8'h00;
			13'h19e1: data_buf = 8'h00;
			13'h19e2: data_buf = 8'h00;
			13'h19e3: data_buf = 8'h81;
			13'h19e4: data_buf = 8'hcd;
			13'h19e5: data_buf = 8'hcd;
			13'h19e6: data_buf = 8'h16;
			13'h19e7: data_buf = 8'h11;
			13'h19e8: data_buf = 8'h8f;
			13'h19e9: data_buf = 8'h15;
			13'h19ea: data_buf = 8'hd5;
			13'h19eb: data_buf = 8'he5;
			13'h19ec: data_buf = 8'hcd;
			13'h19ed: data_buf = 8'he8;
			13'h19ee: data_buf = 8'h16;
			13'h19ef: data_buf = 8'hcd;
			13'h19f0: data_buf = 8'h91;
			13'h19f1: data_buf = 8'h15;
			13'h19f2: data_buf = 8'he1;
			13'h19f3: data_buf = 8'hcd;
			13'h19f4: data_buf = 8'hcd;
			13'h19f5: data_buf = 8'h16;
			13'h19f6: data_buf = 8'h7e;
			13'h19f7: data_buf = 8'h23;
			13'h19f8: data_buf = 8'hcd;
			13'h19f9: data_buf = 8'hda;
			13'h19fa: data_buf = 8'h16;
			13'h19fb: data_buf = 8'h06;
			13'h19fc: data_buf = 8'hf1;
			13'h19fd: data_buf = 8'hc1;
			13'h19fe: data_buf = 8'hd1;
			13'h19ff: data_buf = 8'h3d;
			13'h1a00: data_buf = 8'hc8;
			13'h1a01: data_buf = 8'hd5;
			13'h1a02: data_buf = 8'hc5;
			13'h1a03: data_buf = 8'hf5;
			13'h1a04: data_buf = 8'he5;
			13'h1a05: data_buf = 8'hcd;
			13'h1a06: data_buf = 8'h91;
			13'h1a07: data_buf = 8'h15;
			13'h1a08: data_buf = 8'he1;
			13'h1a09: data_buf = 8'hcd;
			13'h1a0a: data_buf = 8'heb;
			13'h1a0b: data_buf = 8'h16;
			13'h1a0c: data_buf = 8'he5;
			13'h1a0d: data_buf = 8'hcd;
			13'h1a0e: data_buf = 8'h56;
			13'h1a0f: data_buf = 8'h14;
			13'h1a10: data_buf = 8'he1;
			13'h1a11: data_buf = 8'hc3;
			13'h1a12: data_buf = 8'hfc;
			13'h1a13: data_buf = 8'h19;
			13'h1a14: data_buf = 8'hcd;
			13'h1a15: data_buf = 8'h9c;
			13'h1a16: data_buf = 8'h16;
			13'h1a17: data_buf = 8'h21;
			13'h1a18: data_buf = 8'h5e;
			13'h1a19: data_buf = 8'h80;
			13'h1a1a: data_buf = 8'hfa;
			13'h1a1b: data_buf = 8'h75;
			13'h1a1c: data_buf = 8'h1a;
			13'h1a1d: data_buf = 8'h21;
			13'h1a1e: data_buf = 8'h7f;
			13'h1a1f: data_buf = 8'h80;
			13'h1a20: data_buf = 8'hcd;
			13'h1a21: data_buf = 8'hda;
			13'h1a22: data_buf = 8'h16;
			13'h1a23: data_buf = 8'h21;
			13'h1a24: data_buf = 8'h5e;
			13'h1a25: data_buf = 8'h80;
			13'h1a26: data_buf = 8'hc8;
			13'h1a27: data_buf = 8'h86;
			13'h1a28: data_buf = 8'he6;
			13'h1a29: data_buf = 8'h07;
			13'h1a2a: data_buf = 8'h06;
			13'h1a2b: data_buf = 8'h00;
			13'h1a2c: data_buf = 8'h77;
			13'h1a2d: data_buf = 8'h23;
			13'h1a2e: data_buf = 8'h87;
			13'h1a2f: data_buf = 8'h87;
			13'h1a30: data_buf = 8'h4f;
			13'h1a31: data_buf = 8'h09;
			13'h1a32: data_buf = 8'hcd;
			13'h1a33: data_buf = 8'heb;
			13'h1a34: data_buf = 8'h16;
			13'h1a35: data_buf = 8'hcd;
			13'h1a36: data_buf = 8'h91;
			13'h1a37: data_buf = 8'h15;
			13'h1a38: data_buf = 8'h3a;
			13'h1a39: data_buf = 8'h5d;
			13'h1a3a: data_buf = 8'h80;
			13'h1a3b: data_buf = 8'h3c;
			13'h1a3c: data_buf = 8'he6;
			13'h1a3d: data_buf = 8'h03;
			13'h1a3e: data_buf = 8'h06;
			13'h1a3f: data_buf = 8'h00;
			13'h1a40: data_buf = 8'hfe;
			13'h1a41: data_buf = 8'h01;
			13'h1a42: data_buf = 8'h88;
			13'h1a43: data_buf = 8'h32;
			13'h1a44: data_buf = 8'h5d;
			13'h1a45: data_buf = 8'h80;
			13'h1a46: data_buf = 8'h21;
			13'h1a47: data_buf = 8'h79;
			13'h1a48: data_buf = 8'h1a;
			13'h1a49: data_buf = 8'h87;
			13'h1a4a: data_buf = 8'h87;
			13'h1a4b: data_buf = 8'h4f;
			13'h1a4c: data_buf = 8'h09;
			13'h1a4d: data_buf = 8'hcd;
			13'h1a4e: data_buf = 8'h47;
			13'h1a4f: data_buf = 8'h14;
			13'h1a50: data_buf = 8'hcd;
			13'h1a51: data_buf = 8'he8;
			13'h1a52: data_buf = 8'h16;
			13'h1a53: data_buf = 8'h7b;
			13'h1a54: data_buf = 8'h59;
			13'h1a55: data_buf = 8'hee;
			13'h1a56: data_buf = 8'h4f;
			13'h1a57: data_buf = 8'h4f;
			13'h1a58: data_buf = 8'h36;
			13'h1a59: data_buf = 8'h80;
			13'h1a5a: data_buf = 8'h2b;
			13'h1a5b: data_buf = 8'h46;
			13'h1a5c: data_buf = 8'h36;
			13'h1a5d: data_buf = 8'h80;
			13'h1a5e: data_buf = 8'h21;
			13'h1a5f: data_buf = 8'h5c;
			13'h1a60: data_buf = 8'h80;
			13'h1a61: data_buf = 8'h34;
			13'h1a62: data_buf = 8'h7e;
			13'h1a63: data_buf = 8'hd6;
			13'h1a64: data_buf = 8'hab;
			13'h1a65: data_buf = 8'hc2;
			13'h1a66: data_buf = 8'h6c;
			13'h1a67: data_buf = 8'h1a;
			13'h1a68: data_buf = 8'h77;
			13'h1a69: data_buf = 8'h0c;
			13'h1a6a: data_buf = 8'h15;
			13'h1a6b: data_buf = 8'h1c;
			13'h1a6c: data_buf = 8'hcd;
			13'h1a6d: data_buf = 8'ha7;
			13'h1a6e: data_buf = 8'h14;
			13'h1a6f: data_buf = 8'h21;
			13'h1a70: data_buf = 8'h7f;
			13'h1a71: data_buf = 8'h80;
			13'h1a72: data_buf = 8'hc3;
			13'h1a73: data_buf = 8'hf4;
			13'h1a74: data_buf = 8'h16;
			13'h1a75: data_buf = 8'h77;
			13'h1a76: data_buf = 8'h2b;
			13'h1a77: data_buf = 8'h77;
			13'h1a78: data_buf = 8'h2b;
			13'h1a79: data_buf = 8'h77;
			13'h1a7a: data_buf = 8'hc3;
			13'h1a7b: data_buf = 8'h50;
			13'h1a7c: data_buf = 8'h1a;
			13'h1a7d: data_buf = 8'h68;
			13'h1a7e: data_buf = 8'hb1;
			13'h1a7f: data_buf = 8'h46;
			13'h1a80: data_buf = 8'h68;
			13'h1a81: data_buf = 8'h99;
			13'h1a82: data_buf = 8'he9;
			13'h1a83: data_buf = 8'h92;
			13'h1a84: data_buf = 8'h69;
			13'h1a85: data_buf = 8'h10;
			13'h1a86: data_buf = 8'hd1;
			13'h1a87: data_buf = 8'h75;
			13'h1a88: data_buf = 8'h68;
			13'h1a89: data_buf = 8'h21;
			13'h1a8a: data_buf = 8'hd3;
			13'h1a8b: data_buf = 8'h1a;
			13'h1a8c: data_buf = 8'hcd;
			13'h1a8d: data_buf = 8'h47;
			13'h1a8e: data_buf = 8'h14;
			13'h1a8f: data_buf = 8'hcd;
			13'h1a90: data_buf = 8'hcd;
			13'h1a91: data_buf = 8'h16;
			13'h1a92: data_buf = 8'h01;
			13'h1a93: data_buf = 8'h49;
			13'h1a94: data_buf = 8'h83;
			13'h1a95: data_buf = 8'h11;
			13'h1a96: data_buf = 8'hdb;
			13'h1a97: data_buf = 8'h0f;
			13'h1a98: data_buf = 8'hcd;
			13'h1a99: data_buf = 8'hdd;
			13'h1a9a: data_buf = 8'h16;
			13'h1a9b: data_buf = 8'hc1;
			13'h1a9c: data_buf = 8'hd1;
			13'h1a9d: data_buf = 8'hcd;
			13'h1a9e: data_buf = 8'hf2;
			13'h1a9f: data_buf = 8'h15;
			13'h1aa0: data_buf = 8'hcd;
			13'h1aa1: data_buf = 8'hcd;
			13'h1aa2: data_buf = 8'h16;
			13'h1aa3: data_buf = 8'hcd;
			13'h1aa4: data_buf = 8'h6f;
			13'h1aa5: data_buf = 8'h17;
			13'h1aa6: data_buf = 8'hc1;
			13'h1aa7: data_buf = 8'hd1;
			13'h1aa8: data_buf = 8'hcd;
			13'h1aa9: data_buf = 8'h53;
			13'h1aaa: data_buf = 8'h14;
			13'h1aab: data_buf = 8'h21;
			13'h1aac: data_buf = 8'hd7;
			13'h1aad: data_buf = 8'h1a;
			13'h1aae: data_buf = 8'hcd;
			13'h1aaf: data_buf = 8'h4d;
			13'h1ab0: data_buf = 8'h14;
			13'h1ab1: data_buf = 8'hcd;
			13'h1ab2: data_buf = 8'h9c;
			13'h1ab3: data_buf = 8'h16;
			13'h1ab4: data_buf = 8'h37;
			13'h1ab5: data_buf = 8'hf2;
			13'h1ab6: data_buf = 8'hbf;
			13'h1ab7: data_buf = 8'h1a;
			13'h1ab8: data_buf = 8'hcd;
			13'h1ab9: data_buf = 8'h44;
			13'h1aba: data_buf = 8'h14;
			13'h1abb: data_buf = 8'hcd;
			13'h1abc: data_buf = 8'h9c;
			13'h1abd: data_buf = 8'h16;
			13'h1abe: data_buf = 8'hb7;
			13'h1abf: data_buf = 8'hf5;
			13'h1ac0: data_buf = 8'hf4;
			13'h1ac1: data_buf = 8'hc5;
			13'h1ac2: data_buf = 8'h16;
			13'h1ac3: data_buf = 8'h21;
			13'h1ac4: data_buf = 8'hd7;
			13'h1ac5: data_buf = 8'h1a;
			13'h1ac6: data_buf = 8'hcd;
			13'h1ac7: data_buf = 8'h47;
			13'h1ac8: data_buf = 8'h14;
			13'h1ac9: data_buf = 8'hf1;
			13'h1aca: data_buf = 8'hd4;
			13'h1acb: data_buf = 8'hc5;
			13'h1acc: data_buf = 8'h16;
			13'h1acd: data_buf = 8'h21;
			13'h1ace: data_buf = 8'hdb;
			13'h1acf: data_buf = 8'h1a;
			13'h1ad0: data_buf = 8'hc3;
			13'h1ad1: data_buf = 8'he4;
			13'h1ad2: data_buf = 8'h19;
			13'h1ad3: data_buf = 8'hdb;
			13'h1ad4: data_buf = 8'h0f;
			13'h1ad5: data_buf = 8'h49;
			13'h1ad6: data_buf = 8'h81;
			13'h1ad7: data_buf = 8'h00;
			13'h1ad8: data_buf = 8'h00;
			13'h1ad9: data_buf = 8'h00;
			13'h1ada: data_buf = 8'h7f;
			13'h1adb: data_buf = 8'h05;
			13'h1adc: data_buf = 8'hba;
			13'h1add: data_buf = 8'hd7;
			13'h1ade: data_buf = 8'h1e;
			13'h1adf: data_buf = 8'h86;
			13'h1ae0: data_buf = 8'h64;
			13'h1ae1: data_buf = 8'h26;
			13'h1ae2: data_buf = 8'h99;
			13'h1ae3: data_buf = 8'h87;
			13'h1ae4: data_buf = 8'h58;
			13'h1ae5: data_buf = 8'h34;
			13'h1ae6: data_buf = 8'h23;
			13'h1ae7: data_buf = 8'h87;
			13'h1ae8: data_buf = 8'he0;
			13'h1ae9: data_buf = 8'h5d;
			13'h1aea: data_buf = 8'ha5;
			13'h1aeb: data_buf = 8'h86;
			13'h1aec: data_buf = 8'hda;
			13'h1aed: data_buf = 8'h0f;
			13'h1aee: data_buf = 8'h49;
			13'h1aef: data_buf = 8'h83;
			13'h1af0: data_buf = 8'hcd;
			13'h1af1: data_buf = 8'hcd;
			13'h1af2: data_buf = 8'h16;
			13'h1af3: data_buf = 8'hcd;
			13'h1af4: data_buf = 8'h8f;
			13'h1af5: data_buf = 8'h1a;
			13'h1af6: data_buf = 8'hc1;
			13'h1af7: data_buf = 8'he1;
			13'h1af8: data_buf = 8'hcd;
			13'h1af9: data_buf = 8'hcd;
			13'h1afa: data_buf = 8'h16;
			13'h1afb: data_buf = 8'heb;
			13'h1afc: data_buf = 8'hcd;
			13'h1afd: data_buf = 8'hdd;
			13'h1afe: data_buf = 8'h16;
			13'h1aff: data_buf = 8'hcd;
			13'h1b00: data_buf = 8'h89;
			13'h1b01: data_buf = 8'h1a;
			13'h1b02: data_buf = 8'hc3;
			13'h1b03: data_buf = 8'hf0;
			13'h1b04: data_buf = 8'h15;
			13'h1b05: data_buf = 8'hcd;
			13'h1b06: data_buf = 8'h9c;
			13'h1b07: data_buf = 8'h16;
			13'h1b08: data_buf = 8'hfc;
			13'h1b09: data_buf = 8'h30;
			13'h1b0a: data_buf = 8'h19;
			13'h1b0b: data_buf = 8'hfc;
			13'h1b0c: data_buf = 8'hc5;
			13'h1b0d: data_buf = 8'h16;
			13'h1b0e: data_buf = 8'h3a;
			13'h1b0f: data_buf = 8'h2c;
			13'h1b10: data_buf = 8'h81;
			13'h1b11: data_buf = 8'hfe;
			13'h1b12: data_buf = 8'h81;
			13'h1b13: data_buf = 8'hda;
			13'h1b14: data_buf = 8'h22;
			13'h1b15: data_buf = 8'h1b;
			13'h1b16: data_buf = 8'h01;
			13'h1b17: data_buf = 8'h00;
			13'h1b18: data_buf = 8'h81;
			13'h1b19: data_buf = 8'h51;
			13'h1b1a: data_buf = 8'h59;
			13'h1b1b: data_buf = 8'hcd;
			13'h1b1c: data_buf = 8'hf2;
			13'h1b1d: data_buf = 8'h15;
			13'h1b1e: data_buf = 8'h21;
			13'h1b1f: data_buf = 8'h4d;
			13'h1b20: data_buf = 8'h14;
			13'h1b21: data_buf = 8'he5;
			13'h1b22: data_buf = 8'h21;
			13'h1b23: data_buf = 8'h2c;
			13'h1b24: data_buf = 8'h1b;
			13'h1b25: data_buf = 8'hcd;
			13'h1b26: data_buf = 8'he4;
			13'h1b27: data_buf = 8'h19;
			13'h1b28: data_buf = 8'h21;
			13'h1b29: data_buf = 8'hd3;
			13'h1b2a: data_buf = 8'h1a;
			13'h1b2b: data_buf = 8'hc9;
			13'h1b2c: data_buf = 8'h09;
			13'h1b2d: data_buf = 8'h4a;
			13'h1b2e: data_buf = 8'hd7;
			13'h1b2f: data_buf = 8'h3b;
			13'h1b30: data_buf = 8'h78;
			13'h1b31: data_buf = 8'h02;
			13'h1b32: data_buf = 8'h6e;
			13'h1b33: data_buf = 8'h84;
			13'h1b34: data_buf = 8'h7b;
			13'h1b35: data_buf = 8'hfe;
			13'h1b36: data_buf = 8'hc1;
			13'h1b37: data_buf = 8'h2f;
			13'h1b38: data_buf = 8'h7c;
			13'h1b39: data_buf = 8'h74;
			13'h1b3a: data_buf = 8'h31;
			13'h1b3b: data_buf = 8'h9a;
			13'h1b3c: data_buf = 8'h7d;
			13'h1b3d: data_buf = 8'h84;
			13'h1b3e: data_buf = 8'h3d;
			13'h1b3f: data_buf = 8'h5a;
			13'h1b40: data_buf = 8'h7d;
			13'h1b41: data_buf = 8'hc8;
			13'h1b42: data_buf = 8'h7f;
			13'h1b43: data_buf = 8'h91;
			13'h1b44: data_buf = 8'h7e;
			13'h1b45: data_buf = 8'he4;
			13'h1b46: data_buf = 8'hbb;
			13'h1b47: data_buf = 8'h4c;
			13'h1b48: data_buf = 8'h7e;
			13'h1b49: data_buf = 8'h6c;
			13'h1b4a: data_buf = 8'haa;
			13'h1b4b: data_buf = 8'haa;
			13'h1b4c: data_buf = 8'h7f;
			13'h1b4d: data_buf = 8'h00;
			13'h1b4e: data_buf = 8'h00;
			13'h1b4f: data_buf = 8'h00;
			13'h1b50: data_buf = 8'h81;
			13'h1b51: data_buf = 8'hc9;
			13'h1b52: data_buf = 8'hd7;
			13'h1b53: data_buf = 8'hc9;
			13'h1b54: data_buf = 8'h3e;
			13'h1b55: data_buf = 8'h0c;
			13'h1b56: data_buf = 8'hc3;
			13'h1b57: data_buf = 8'h8a;
			13'h1b58: data_buf = 8'h1c;
			13'h1b59: data_buf = 8'hcd;
			13'h1b5a: data_buf = 8'h1b;
			13'h1b5b: data_buf = 8'h14;
			13'h1b5c: data_buf = 8'h7b;
			13'h1b5d: data_buf = 8'h32;
			13'h1b5e: data_buf = 8'h87;
			13'h1b5f: data_buf = 8'h80;
			13'h1b60: data_buf = 8'hc9;
			13'h1b61: data_buf = 8'hcd;
			13'h1b62: data_buf = 8'hba;
			13'h1b63: data_buf = 8'h0c;
			13'h1b64: data_buf = 8'hcd;
			13'h1b65: data_buf = 8'hff;
			13'h1b66: data_buf = 8'h08;
			13'h1b67: data_buf = 8'hed;
			13'h1b68: data_buf = 8'h53;
			13'h1b69: data_buf = 8'h8b;
			13'h1b6a: data_buf = 8'h80;
			13'h1b6b: data_buf = 8'hed;
			13'h1b6c: data_buf = 8'h53;
			13'h1b6d: data_buf = 8'h8d;
			13'h1b6e: data_buf = 8'h80;
			13'h1b6f: data_buf = 8'hc9;
			13'h1b70: data_buf = 8'hcd;
			13'h1b71: data_buf = 8'hff;
			13'h1b72: data_buf = 8'h08;
			13'h1b73: data_buf = 8'hd5;
			13'h1b74: data_buf = 8'he1;
			13'h1b75: data_buf = 8'h46;
			13'h1b76: data_buf = 8'h23;
			13'h1b77: data_buf = 8'h7e;
			13'h1b78: data_buf = 8'hc3;
			13'h1b79: data_buf = 8'h75;
			13'h1b7a: data_buf = 8'h10;
			13'h1b7b: data_buf = 8'hcd;
			13'h1b7c: data_buf = 8'hba;
			13'h1b7d: data_buf = 8'h0c;
			13'h1b7e: data_buf = 8'hcd;
			13'h1b7f: data_buf = 8'hff;
			13'h1b80: data_buf = 8'h08;
			13'h1b81: data_buf = 8'hd5;
			13'h1b82: data_buf = 8'hcd;
			13'h1b83: data_buf = 8'hc3;
			13'h1b84: data_buf = 8'h06;
			13'h1b85: data_buf = 8'h2c;
			13'h1b86: data_buf = 8'hcd;
			13'h1b87: data_buf = 8'hba;
			13'h1b88: data_buf = 8'h0c;
			13'h1b89: data_buf = 8'hcd;
			13'h1b8a: data_buf = 8'hff;
			13'h1b8b: data_buf = 8'h08;
			13'h1b8c: data_buf = 8'he3;
			13'h1b8d: data_buf = 8'h73;
			13'h1b8e: data_buf = 8'h23;
			13'h1b8f: data_buf = 8'h72;
			13'h1b90: data_buf = 8'he1;
			13'h1b91: data_buf = 8'hc9;
			13'h1b92: data_buf = 8'hcd;
			13'h1b93: data_buf = 8'hbd;
			13'h1b94: data_buf = 8'h0c;
			13'h1b95: data_buf = 8'hcd;
			13'h1b96: data_buf = 8'hff;
			13'h1b97: data_buf = 8'h08;
			13'h1b98: data_buf = 8'hc5;
			13'h1b99: data_buf = 8'h21;
			13'h1b9a: data_buf = 8'h2e;
			13'h1b9b: data_buf = 8'h81;
			13'h1b9c: data_buf = 8'h7a;
			13'h1b9d: data_buf = 8'hfe;
			13'h1b9e: data_buf = 8'h00;
			13'h1b9f: data_buf = 8'h28;
			13'h1ba0: data_buf = 8'h0c;
			13'h1ba1: data_buf = 8'hcd;
			13'h1ba2: data_buf = 8'hca;
			13'h1ba3: data_buf = 8'h1b;
			13'h1ba4: data_buf = 8'h78;
			13'h1ba5: data_buf = 8'hfe;
			13'h1ba6: data_buf = 8'h30;
			13'h1ba7: data_buf = 8'h28;
			13'h1ba8: data_buf = 8'h02;
			13'h1ba9: data_buf = 8'h70;
			13'h1baa: data_buf = 8'h23;
			13'h1bab: data_buf = 8'h71;
			13'h1bac: data_buf = 8'h23;
			13'h1bad: data_buf = 8'h7b;
			13'h1bae: data_buf = 8'hcd;
			13'h1baf: data_buf = 8'hca;
			13'h1bb0: data_buf = 8'h1b;
			13'h1bb1: data_buf = 8'h7a;
			13'h1bb2: data_buf = 8'hfe;
			13'h1bb3: data_buf = 8'h00;
			13'h1bb4: data_buf = 8'h20;
			13'h1bb5: data_buf = 8'h05;
			13'h1bb6: data_buf = 8'h78;
			13'h1bb7: data_buf = 8'hfe;
			13'h1bb8: data_buf = 8'h30;
			13'h1bb9: data_buf = 8'h28;
			13'h1bba: data_buf = 8'h02;
			13'h1bbb: data_buf = 8'h70;
			13'h1bbc: data_buf = 8'h23;
			13'h1bbd: data_buf = 8'h71;
			13'h1bbe: data_buf = 8'h23;
			13'h1bbf: data_buf = 8'haf;
			13'h1bc0: data_buf = 8'h77;
			13'h1bc1: data_buf = 8'h23;
			13'h1bc2: data_buf = 8'h77;
			13'h1bc3: data_buf = 8'hc1;
			13'h1bc4: data_buf = 8'h21;
			13'h1bc5: data_buf = 8'h2e;
			13'h1bc6: data_buf = 8'h81;
			13'h1bc7: data_buf = 8'hc3;
			13'h1bc8: data_buf = 8'h23;
			13'h1bc9: data_buf = 8'h11;
			13'h1bca: data_buf = 8'h47;
			13'h1bcb: data_buf = 8'he6;
			13'h1bcc: data_buf = 8'h0f;
			13'h1bcd: data_buf = 8'hfe;
			13'h1bce: data_buf = 8'h0a;
			13'h1bcf: data_buf = 8'h38;
			13'h1bd0: data_buf = 8'h02;
			13'h1bd1: data_buf = 8'hc6;
			13'h1bd2: data_buf = 8'h07;
			13'h1bd3: data_buf = 8'hc6;
			13'h1bd4: data_buf = 8'h30;
			13'h1bd5: data_buf = 8'h4f;
			13'h1bd6: data_buf = 8'h78;
			13'h1bd7: data_buf = 8'h0f;
			13'h1bd8: data_buf = 8'h0f;
			13'h1bd9: data_buf = 8'h0f;
			13'h1bda: data_buf = 8'h0f;
			13'h1bdb: data_buf = 8'he6;
			13'h1bdc: data_buf = 8'h0f;
			13'h1bdd: data_buf = 8'hfe;
			13'h1bde: data_buf = 8'h0a;
			13'h1bdf: data_buf = 8'h38;
			13'h1be0: data_buf = 8'h02;
			13'h1be1: data_buf = 8'hc6;
			13'h1be2: data_buf = 8'h07;
			13'h1be3: data_buf = 8'hc6;
			13'h1be4: data_buf = 8'h30;
			13'h1be5: data_buf = 8'h47;
			13'h1be6: data_buf = 8'hc9;
			13'h1be7: data_buf = 8'heb;
			13'h1be8: data_buf = 8'h21;
			13'h1be9: data_buf = 8'h00;
			13'h1bea: data_buf = 8'h00;
			13'h1beb: data_buf = 8'hcd;
			13'h1bec: data_buf = 8'h00;
			13'h1bed: data_buf = 8'h1c;
			13'h1bee: data_buf = 8'hda;
			13'h1bef: data_buf = 8'h20;
			13'h1bf0: data_buf = 8'h1c;
			13'h1bf1: data_buf = 8'h18;
			13'h1bf2: data_buf = 8'h05;
			13'h1bf3: data_buf = 8'hcd;
			13'h1bf4: data_buf = 8'h00;
			13'h1bf5: data_buf = 8'h1c;
			13'h1bf6: data_buf = 8'h38;
			13'h1bf7: data_buf = 8'h1f;
			13'h1bf8: data_buf = 8'h29;
			13'h1bf9: data_buf = 8'h29;
			13'h1bfa: data_buf = 8'h29;
			13'h1bfb: data_buf = 8'h29;
			13'h1bfc: data_buf = 8'hb5;
			13'h1bfd: data_buf = 8'h6f;
			13'h1bfe: data_buf = 8'h18;
			13'h1bff: data_buf = 8'hf3;
			13'h1c00: data_buf = 8'h13;
			13'h1c01: data_buf = 8'h1a;
			13'h1c02: data_buf = 8'hfe;
			13'h1c03: data_buf = 8'h20;
			13'h1c04: data_buf = 8'hca;
			13'h1c05: data_buf = 8'h00;
			13'h1c06: data_buf = 8'h1c;
			13'h1c07: data_buf = 8'hd6;
			13'h1c08: data_buf = 8'h30;
			13'h1c09: data_buf = 8'hd8;
			13'h1c0a: data_buf = 8'hfe;
			13'h1c0b: data_buf = 8'h0a;
			13'h1c0c: data_buf = 8'h38;
			13'h1c0d: data_buf = 8'h05;
			13'h1c0e: data_buf = 8'hd6;
			13'h1c0f: data_buf = 8'h07;
			13'h1c10: data_buf = 8'hfe;
			13'h1c11: data_buf = 8'h0a;
			13'h1c12: data_buf = 8'hd8;
			13'h1c13: data_buf = 8'hfe;
			13'h1c14: data_buf = 8'h10;
			13'h1c15: data_buf = 8'h3f;
			13'h1c16: data_buf = 8'hc9;
			13'h1c17: data_buf = 8'heb;
			13'h1c18: data_buf = 8'h7a;
			13'h1c19: data_buf = 8'h4b;
			13'h1c1a: data_buf = 8'he5;
			13'h1c1b: data_buf = 8'hcd;
			13'h1c1c: data_buf = 8'h74;
			13'h1c1d: data_buf = 8'h10;
			13'h1c1e: data_buf = 8'he1;
			13'h1c1f: data_buf = 8'hc9;
			13'h1c20: data_buf = 8'h1e;
			13'h1c21: data_buf = 8'h26;
			13'h1c22: data_buf = 8'hc3;
			13'h1c23: data_buf = 8'h09;
			13'h1c24: data_buf = 8'h04;
			13'h1c25: data_buf = 8'hcd;
			13'h1c26: data_buf = 8'hbd;
			13'h1c27: data_buf = 8'h0c;
			13'h1c28: data_buf = 8'hcd;
			13'h1c29: data_buf = 8'hff;
			13'h1c2a: data_buf = 8'h08;
			13'h1c2b: data_buf = 8'hc5;
			13'h1c2c: data_buf = 8'h21;
			13'h1c2d: data_buf = 8'h2e;
			13'h1c2e: data_buf = 8'h81;
			13'h1c2f: data_buf = 8'h06;
			13'h1c30: data_buf = 8'h11;
			13'h1c31: data_buf = 8'h05;
			13'h1c32: data_buf = 8'h78;
			13'h1c33: data_buf = 8'hfe;
			13'h1c34: data_buf = 8'h01;
			13'h1c35: data_buf = 8'h28;
			13'h1c36: data_buf = 8'h08;
			13'h1c37: data_buf = 8'hcb;
			13'h1c38: data_buf = 8'h13;
			13'h1c39: data_buf = 8'hcb;
			13'h1c3a: data_buf = 8'h12;
			13'h1c3b: data_buf = 8'h30;
			13'h1c3c: data_buf = 8'hf4;
			13'h1c3d: data_buf = 8'h18;
			13'h1c3e: data_buf = 8'h04;
			13'h1c3f: data_buf = 8'hcb;
			13'h1c40: data_buf = 8'h13;
			13'h1c41: data_buf = 8'hcb;
			13'h1c42: data_buf = 8'h12;
			13'h1c43: data_buf = 8'h3e;
			13'h1c44: data_buf = 8'h30;
			13'h1c45: data_buf = 8'hce;
			13'h1c46: data_buf = 8'h00;
			13'h1c47: data_buf = 8'h77;
			13'h1c48: data_buf = 8'h23;
			13'h1c49: data_buf = 8'h05;
			13'h1c4a: data_buf = 8'h20;
			13'h1c4b: data_buf = 8'hf3;
			13'h1c4c: data_buf = 8'haf;
			13'h1c4d: data_buf = 8'h77;
			13'h1c4e: data_buf = 8'h23;
			13'h1c4f: data_buf = 8'h77;
			13'h1c50: data_buf = 8'hc1;
			13'h1c51: data_buf = 8'h21;
			13'h1c52: data_buf = 8'h2e;
			13'h1c53: data_buf = 8'h81;
			13'h1c54: data_buf = 8'hc3;
			13'h1c55: data_buf = 8'h23;
			13'h1c56: data_buf = 8'h11;
			13'h1c57: data_buf = 8'heb;
			13'h1c58: data_buf = 8'h21;
			13'h1c59: data_buf = 8'h00;
			13'h1c5a: data_buf = 8'h00;
			13'h1c5b: data_buf = 8'hcd;
			13'h1c5c: data_buf = 8'h74;
			13'h1c5d: data_buf = 8'h1c;
			13'h1c5e: data_buf = 8'hda;
			13'h1c5f: data_buf = 8'h82;
			13'h1c60: data_buf = 8'h1c;
			13'h1c61: data_buf = 8'hd6;
			13'h1c62: data_buf = 8'h30;
			13'h1c63: data_buf = 8'h29;
			13'h1c64: data_buf = 8'hb5;
			13'h1c65: data_buf = 8'h6f;
			13'h1c66: data_buf = 8'hcd;
			13'h1c67: data_buf = 8'h74;
			13'h1c68: data_buf = 8'h1c;
			13'h1c69: data_buf = 8'h30;
			13'h1c6a: data_buf = 8'hf6;
			13'h1c6b: data_buf = 8'heb;
			13'h1c6c: data_buf = 8'h7a;
			13'h1c6d: data_buf = 8'h4b;
			13'h1c6e: data_buf = 8'he5;
			13'h1c6f: data_buf = 8'hcd;
			13'h1c70: data_buf = 8'h74;
			13'h1c71: data_buf = 8'h10;
			13'h1c72: data_buf = 8'he1;
			13'h1c73: data_buf = 8'hc9;
			13'h1c74: data_buf = 8'h13;
			13'h1c75: data_buf = 8'h1a;
			13'h1c76: data_buf = 8'hfe;
			13'h1c77: data_buf = 8'h20;
			13'h1c78: data_buf = 8'hca;
			13'h1c79: data_buf = 8'h74;
			13'h1c7a: data_buf = 8'h1c;
			13'h1c7b: data_buf = 8'hfe;
			13'h1c7c: data_buf = 8'h30;
			13'h1c7d: data_buf = 8'hd8;
			13'h1c7e: data_buf = 8'hfe;
			13'h1c7f: data_buf = 8'h32;
			13'h1c80: data_buf = 8'h3f;
			13'h1c81: data_buf = 8'hc9;
			13'h1c82: data_buf = 8'h1e;
			13'h1c83: data_buf = 8'h28;
			13'h1c84: data_buf = 8'hc3;
			13'h1c85: data_buf = 8'h09;
			13'h1c86: data_buf = 8'h04;
			13'h1c87: data_buf = 8'hc3;
			13'h1c88: data_buf = 8'h4e;
			13'h1c89: data_buf = 8'h00;
			13'h1c8a: data_buf = 8'hc3;
			13'h1c8b: data_buf = 8'h08;
			13'h1c8c: data_buf = 8'h00;
			13'h1c8d: data_buf = 8'hc3;
			13'h1c8e: data_buf = 8'h00;
			13'h1c8f: data_buf = 8'h00;
			13'h1c90: data_buf = 8'h3e;
			13'h1c91: data_buf = 8'h00;
			13'h1c92: data_buf = 8'h32;
			13'h1c93: data_buf = 8'h92;
			13'h1c94: data_buf = 8'h80;
			13'h1c95: data_buf = 8'hc3;
			13'h1c96: data_buf = 8'h55;
			13'h1c97: data_buf = 8'h00;
			13'h1c98: data_buf = 8'hf5;
			13'h1c99: data_buf = 8'ha0;
			13'h1c9a: data_buf = 8'hc1;
			13'h1c9b: data_buf = 8'hb8;
			13'h1c9c: data_buf = 8'h3e;
			13'h1c9d: data_buf = 8'h00;
			13'h1c9e: data_buf = 8'hc9;
			13'h1c9f: data_buf = 8'hcd;
			13'h1ca0: data_buf = 8'hce;
			13'h1ca1: data_buf = 8'h06;
			13'h1ca2: data_buf = 8'hc3;
			13'h1ca3: data_buf = 8'hf5;
			13'h1ca4: data_buf = 8'h0a;

			default:  data_buf = 8'hFF;
		endcase
	end
end

assign data = (ce & oe) ? data_buf : 8'hzz;

endmodule